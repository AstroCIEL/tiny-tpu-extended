// ===== MLP量化参数（SystemVerilog参数定义）=====
// 第1层权重 (int8)
logic signed [7:0] layer1_weight [0:63][0:255] = '{
    '{4, 5, -5, 27, 45, 77, 55, 17, 10, 58, 83, 79, 85, 47, 1, -4, -20, -2, -9, 30, 16, 35, 47, 20, 20, 17, 2, -8, 15, 35, 1, -13, 6, -3, 14, 20, 11, 18, 12, 5, -7, -4, 3, 8, 4, 3, -16, 8, -24, -19, -1, -24, -28, -13, -11, -23, -12, -4, 6, 7, 0, -2, -3, -4, -24, -17, 3, -23, -29, -9, -10, -11, -2, -4, -4, -1, -3, -22, -12, -3, -24, 8, 9, -2, -7, 4, -8, 7, 4, -12, -11, -1, -9, -11, -26, -30, -10, -4, 8, 20, 4, -7, -5, -14, -19, -18, -15, -4, 3, 9, 0, -52, -6, -11, -7, 4, 6, 3, -16, -8, -3, 0, -9, 2, 15, 30, 8, -26, -40, 21, -7, 9, 15, 16, 14, 24, 17, 13, 2, 13, 14, -3, 9, 40, -2, 31, -6, -1, 10, 16, 31, 24, 20, 9, 5, 7, 1, 0, 29, 36, -39, -8, -17, -18, -1, -1, -1, -4, 8, 6, 7, -7, -8, 3, 14, 13, -31, -11, -15, -15, 7, 13, 13, 0, 28, 21, 21, 6, 7, 21, 10, 51, 28, 28, -2, 1, 12, 14, 8, 16, 14, 14, 17, 6, -4, 13, -1, 17, 11, -18, -26, -8, 8, 15, -4, -2, -5, -13, -7, 2, 8, 7, -4, -15, -15, -39, -41, -2, -2, -6, -19, -20, -21, -28, -32, -18, -17, -24, -22, 32, -4, 17, 35, 41, 6, -15, 7, 17, 2, 3, -1, -12, 0, -2, -45, 9},
    '{0, -3, -11, -17, -18, -20, -23, 13, 33, -12, -14, -1, -42, -25, -14, -3, 9, -10, 0, -4, 9, -19, -22, -2, 8, 2, 10, 20, 2, -25, -39, -34, -22, -31, 20, 25, 20, 15, 5, -8, -2, 8, 3, 19, 22, 12, 15, 1, 17, -9, -10, 14, 8, 14, -8, -25, -23, 3, 15, 31, 8, -2, 6, 23, -28, 1, -1, 11, 1, 6, 2, -27, -13, 17, 14, 17, 7, -14, -16, 11, -14, -11, 5, 3, 11, 19, 10, -15, -3, 11, -4, -14, 4, -26, -9, -3, 41, -5, -6, 7, 5, 16, 6, -10, 1, 10, -12, -24, -15, -44, -42, -4, 67, -3, 9, 12, 15, -9, -12, -40, -4, 13, -8, -9, 0, -12, -30, -12, 41, 7, 9, 8, 10, 4, -19, -27, 7, 16, -2, -5, 15, 27, -12, 1, -1, -8, -9, 0, 16, 12, -19, -35, 17, 9, 5, 3, 10, 14, -7, -2, 21, 12, -2, 1, 3, 5, -25, -35, 24, 15, 5, 13, 9, 1, 8, -42, -26, 6, -7, 7, 7, 2, -18, -18, 22, 20, 8, 11, 6, 7, 17, -45, -48, -44, -25, -11, -7, -6, -7, 5, 27, 23, 19, 16, 20, -2, 14, -4, -39, -57, -35, -23, -46, -16, -9, 0, 16, 20, 19, 16, -6, -25, 9, 30, -15, 2, 1, -42, -51, -21, 1, 12, 11, 11, 11, -2, -8, -18, -49, -21, 4, 6, 7, -25, 17, 29, 10, 18, 25, 18, 16, 8, 18, 18, -40, -9},
    '{-3, 0, 9, -11, -28, -37, 3, 16, -31, -41, -46, -46, -32, -40, -24, 1, -31, -20, 25, -5, 8, 4, 8, 13, 19, -6, -14, -2, 7, -31, -36, 1, -39, -34, -26, -19, 10, 20, 15, -6, 6, 16, 10, 1, 7, -4, 4, 22, -49, -42, 11, 2, 2, -8, -12, 1, 6, 16, 3, -7, 2, 12, -14, -10, 29, 20, 13, 3, -10, -8, -12, 3, 7, 22, 11, -2, 9, 28, 28, -14, 14, 26, -22, -21, -9, 6, 2, 3, 4, 18, 12, 12, 8, 15, 13, -44, -11, -7, -25, -10, 5, 16, -5, 14, 1, -3, -6, -16, -11, 0, -7, -52, -24, -3, -2, 21, 18, 16, 12, 10, -22, -25, -3, -1, 0, -1, 8, -39, -16, -18, 5, 17, 28, 15, 11, -1, -20, -10, 14, 6, 2, 4, 28, -13, 11, 6, 4, -2, -1, 6, 27, -7, -20, 13, 12, 7, 15, 17, 16, -19, -19, 12, 13, 7, 7, 14, 25, 5, -10, 8, -5, 2, 15, 1, -41, -49, 11, 27, 14, 1, 10, 7, 20, 24, 7, -1, -4, 1, 26, -5, -46, -25, 13, 21, 17, 1, 0, -8, 8, 9, -3, -4, 1, 3, 28, 9, -25, 21, 15, 54, 12, -8, -2, -7, 8, 7, 10, 5, 10, 10, 15, 0, -32, -3, -15, 14, 2, 9, -3, -4, 13, 11, 16, -3, -5, -12, -5, -1, -37, -35, 4, -4, 32, 32, -20, -47, -19, -16, -30, -22, -14, -46, -19, -14, -17, 0},
    '{-2, -3, -30, 11, 20, 35, 13, 22, 47, 34, 24, 15, 11, 3, 17, 1, 25, -6, -52, -36, -17, 14, 22, 14, 9, 4, -10, -30, -15, 13, -9, -16, 28, 6, 12, 19, 7, 4, 9, 17, 2, -1, -3, -8, -7, -2, -2, -22, -37, -11, 7, -3, -9, -1, 2, -4, -3, -1, 6, 0, 2, -1, -6, -35, -38, -6, 4, -9, -16, -10, -6, 9, 4, -6, -6, -5, -3, -3, -14, 6, -31, 18, -1, 3, -11, -10, -8, 15, 16, 16, 3, -3, -2, 12, -22, 9, -13, 5, 7, 18, -4, -10, 0, -2, 5, -7, -16, 6, 14, 13, -6, -20, -26, -2, -5, 2, -10, -10, -20, -11, -5, -7, -13, 2, 20, 9, 8, 4, -58, 14, -12, -8, -9, -12, -11, 10, 11, 3, -2, 4, 5, -17, -10, 45, -1, 16, -4, 6, 4, 16, 20, 21, 21, 7, 2, 7, 1, -15, -5, 42, -49, -11, -2, -1, 6, 13, 0, 7, 8, 3, 10, 5, -3, -1, 7, 24, -41, -4, -1, 4, 6, 5, 4, 3, 22, 21, 17, 11, 3, 12, 9, 38, 25, 37, 17, 18, 20, 6, 4, -6, 1, 4, 11, 10, 8, 19, 7, -9, 20, -20, -6, 15, 17, 8, 10, 7, -1, -8, 7, 13, 26, 19, 2, -11, -18, -44, -33, -2, -9, -15, -28, -23, -7, -13, -15, -13, -9, -20, -15, 29, 3, 1, 19, 27, 11, -9, -6, -12, -7, -16, -21, -26, -13, -32, -54, 9},
    '{-3, 2, -34, -14, 6, 4, -30, 9, 17, 7, -5, -39, -33, -39, 3, -1, -1, -32, -50, -18, -8, -5, -5, 1, 1, 13, -1, -27, -25, -56, -34, -17, -23, -52, -15, 27, 2, 1, 5, 1, 10, 19, 11, 1, -4, -16, -1, -7, 18, 4, 1, 14, 5, 16, 6, 4, 8, 17, 24, 11, 5, 14, 1, 10, -19, 11, -27, -2, 1, 9, 6, 2, 2, 18, 23, 20, 8, 6, -30, 6, -37, -30, -41, -10, -15, -17, -17, -31, -38, 15, 30, 10, 0, -4, -79, -22, -50, -62, -57, -52, -54, -41, -28, -34, -44, 14, 16, 14, -2, -25, -38, -8, -44, -26, -54, -40, -31, -8, 5, 2, -9, -3, -6, -4, -18, -16, 31, 25, -28, 14, -2, 17, 21, 14, 2, -10, -10, 5, 2, -9, -24, 3, 29, 40, 3, -5, 8, 19, 13, 9, -2, -20, -5, 10, 5, 0, 1, -10, 9, 23, 12, -5, -5, 5, 12, 22, 11, 9, 16, 11, 19, 12, 2, -14, 37, 36, -37, -2, -5, 2, 0, 3, 10, 19, 7, 8, 6, 10, 0, -7, 23, 20, -5, 0, -4, -4, -11, -14, 3, 1, -8, 8, 9, 19, 21, 5, 7, -25, 24, -32, -15, 1, -12, -15, 3, -2, -22, -14, -21, -13, 9, -5, -11, -20, 20, -4, 16, -11, -12, 4, 21, 11, -20, -7, -40, -35, 18, -9, 14, 19, 2, 17, -25, -35, 29, 67, 22, -2, 15, 14, -32, -36, -7, -32, 7, 10},
    '{2, 3, 3, -3, 13, 0, -26, -29, -33, -19, -23, -46, -40, -34, 15, -4, -24, -26, 21, 18, 20, 11, 8, -5, 5, -4, -12, -10, -12, -22, 4, -8, -26, 5, -22, 2, 6, 19, 29, 4, 11, 31, 26, 8, 2, -9, 3, -5, 2, 6, 10, 6, -1, -1, 3, 2, 5, 19, 7, 4, -6, -5, 10, 37, 16, -5, 24, 20, 14, 11, 2, -10, 3, 8, 2, 1, 2, 10, 16, 39, -8, -3, -1, 4, 5, 5, -4, -3, -15, 5, 7, 6, 23, 33, 25, 29, -31, 12, 9, -16, -17, -3, 11, 4, -13, -1, 7, -11, -14, -16, -20, 12, -22, 18, 0, 2, -13, 3, 22, 15, -7, -5, 4, -5, -24, -45, -54, -17, 38, 5, 8, 2, 3, 10, 5, 7, 12, 12, -3, -14, -21, -5, 29, 31, 48, 34, 15, -7, -19, -16, -31, -9, 0, 9, 13, 15, 28, 27, 53, 34, -4, 37, 32, 8, -12, -19, -31, -37, -22, 1, 9, 3, 2, -2, -1, -28, 12, 39, 22, 11, -6, 7, 4, -4, -15, 2, 1, -10, 7, 18, 8, 20, 4, 25, -2, 1, 6, 0, 22, 15, -2, -9, -1, 2, 25, 36, 6, 31, 32, 61, 4, -11, 2, 15, 21, 19, 11, 6, 9, 6, 15, 20, -11, -2, -19, 27, -33, -13, -6, 0, 5, 27, 10, 7, 13, -1, 2, 9, 15, 0, 0, 0, -61, -49, -55, -69, -16, -39, -51, -6, 2, 0, -34, -16, 5, 9},
    '{-1, -1, 14, 8, -22, -36, -42, 9, 55, 33, 72, 104, 127, 53, 18, 3, 27, 54, 39, -33, -58, -73, -83, -13, 3, 11, 37, 29, -7, -14, -35, -36, 43, 43, -31, -43, -44, -31, -34, 8, 9, 0, 12, 1, -27, -46, -44, -45, 5, -1, -53, -32, -35, -35, -21, -2, 15, 8, 2, -21, -24, -34, -27, -52, -29, -33, -26, -22, -38, -29, -6, 19, 28, 9, -11, -16, 12, -14, -32, -7, -19, -31, -39, -23, -28, -3, 5, 25, 39, -28, -51, -23, -7, 1, -17, 20, -22, -21, -51, -30, -3, 11, 11, 22, 23, -21, -12, -21, -6, -10, -39, -5, -6, -19, -35, -22, -4, 7, -4, 7, 13, -3, 3, -15, -13, -24, -46, -56, -7, -31, -24, -43, -15, 12, 8, 21, 2, -2, -10, 2, -7, -42, -38, -28, 17, -14, -22, -36, 9, 19, 20, 3, 3, -19, -26, -16, -21, -12, -4, -46, -5, 10, -10, -18, -3, 17, 1, 11, 17, -32, -23, 0, 4, 30, 9, -19, -22, 0, -10, 17, -5, -10, 0, 12, 17, -17, -5, 13, 19, 35, 31, -7, 4, -10, -14, -16, -6, -11, -9, 8, 8, 0, 6, 12, 25, 13, 22, 9, 4, -5, -20, -47, -39, -19, -18, 3, 0, 15, 12, -6, 0, 2, 8, 29, 4, -1, -27, -35, -24, -26, -15, -21, -10, 8, -4, -36, -34, -2, 21, 20, -2, 3, 6, -4, 15, 10, 11, 16, 28, 8, -10, -22, -20, -30, -7, -14},
    '{3, -2, -10, 4, 17, -10, -36, -30, 5, -16, -37, -73, -75, -17, 10, -4, 8, -9, -14, -1, -6, 7, 18, 15, 1, -8, -8, 0, -3, -39, -9, 6, -4, -14, 1, -29, -31, -13, -22, -8, -8, 1, 0, -7, -15, -9, -2, -29, -10, -18, -16, -41, -46, -26, -19, -22, -9, -17, -23, -5, 0, -3, 3, 15, -47, -19, -12, -16, -23, -11, -18, -13, 3, 6, 7, 13, 17, 16, 19, 18, -30, 5, 10, 1, -8, -15, -12, -2, 17, 22, 21, 25, 15, 14, 29, 4, -34, -31, 5, 6, 5, 13, 12, -1, 8, -6, -32, -19, -13, -5, 27, 41, -23, -13, -18, 8, 17, 19, 9, 9, 16, 22, -11, -23, -37, -39, -1, 40, -9, -6, -5, 9, 8, 13, 2, 10, 19, 22, 3, -22, -29, -15, 4, 40, -9, 10, 3, 11, -2, 1, 12, 11, 5, -15, -25, -13, 2, -2, 10, 42, -67, 9, 2, 1, -2, 8, 13, 12, 4, -12, -19, 2, -7, -11, -1, 0, -52, -17, -12, -23, -24, -15, -5, 0, 6, 12, 21, 8, -20, -2, 52, 17, -43, -42, -11, -8, -25, -13, -4, 0, 9, 12, 19, 14, -18, -6, 46, -12, 13, -24, -24, -21, -27, -5, -3, 10, 3, 7, 15, 20, -7, 7, 42, 16, 7, -17, -77, -69, -47, -25, -14, -5, 1, 3, 32, 26, 46, 40, 50, 32, 1, -4, -10, -24, -20, -50, -14, 16, -4, 6, -16, -1, 0, 7, 37, 9},
    '{-4, -1, -15, 38, 30, 39, 37, -1, -9, 3, 52, 57, 89, 59, -14, -1, -27, -29, 0, 47, 24, 23, 36, 12, 24, 16, 7, 2, 24, 35, -1, -1, -16, -26, 10, 21, 20, 14, 10, 10, 4, 4, -1, 9, 10, 11, 1, 9, 13, 7, 25, -2, 7, 9, -3, -6, -1, 17, 11, -3, -8, 3, 13, 9, -18, 2, 33, 13, 6, 10, 1, -13, -9, 3, 6, 0, -12, -16, -6, 1, -5, -27, 10, 1, -5, 6, -14, -23, -16, -18, -17, -1, -1, -6, -17, 8, -16, -32, -8, 3, 9, 9, -13, -9, -2, -5, -24, -13, 1, 1, -7, -23, -14, -9, -16, -2, 5, 5, 6, 6, 13, 5, -15, -4, 15, 27, 9, -21, -7, 15, -6, 15, 11, 9, 9, 22, 22, 7, -1, 15, 21, 15, -7, -1, 11, 24, -8, 16, 33, 24, 14, 13, 20, 9, 9, 12, 20, 3, 14, 22, -4, 7, 14, -1, 4, 1, -12, -2, -3, 3, 9, -2, 2, 6, 25, 19, -34, -19, -5, -12, -13, -10, -13, -26, 0, 6, -6, -15, -18, -26, -28, 5, -29, -45, -29, -10, -4, 6, -1, 6, 13, 5, -8, -10, -11, -33, -24, 5, 28, -31, -31, 4, 21, 14, 1, 15, 7, -8, -13, -4, -7, -23, -27, -15, 26, -6, -30, -11, -27, -21, -4, -9, 6, -11, -7, -29, -19, -22, -22, 38, 2, -2, -41, -31, -23, -21, -9, -28, -27, -12, -5, -47, -47, -35, -46, 11},
    '{2, -3, 1, 22, 16, 15, 12, 20, 50, 70, 69, 22, -30, 13, 23, -1, 1, -2, -32, -20, -15, -32, -12, -35, -37, -12, 15, -7, -20, -19, 1, -2, 5, -1, 32, -16, -13, 2, -13, -7, 0, 7, 2, 3, 0, -1, 8, 8, 12, 29, 24, -19, -9, 7, -3, -5, -7, 4, -7, 1, 4, 2, -1, 18, 32, 0, -13, -21, -8, 7, 11, 11, 1, 4, 9, 8, 6, 14, -24, -11, 40, -8, 12, 20, 5, 17, 22, 28, 13, 22, 18, 6, 8, 27, -13, -13, 25, 15, 17, 26, 5, 11, 1, -34, -47, -1, -3, -3, 5, -20, -31, 15, 35, 7, -25, -4, -3, -19, -37, -58, -16, -3, -12, -21, -21, -36, -36, -12, 20, -19, -61, -43, -27, -42, -29, -7, 7, 0, 4, -6, 6, 1, -13, 20, -17, -31, -55, -25, -6, -1, -16, -11, 1, -3, -2, 0, 17, 14, 10, 7, -2, 10, 3, 7, 27, 10, -9, -10, 2, -8, -10, 0, -3, 5, 13, 9, 1, 35, 33, 22, 18, 13, 6, 3, 6, -2, -14, 12, 5, 5, 7, 15, 10, 5, 17, 8, 1, 13, 9, 16, 16, 17, 15, 15, 15, 23, 24, 7, 36, -11, 14, 28, -3, -5, -5, -2, 2, 2, 3, -7, 1, 20, 11, -7, 6, 13, 25, 2, 17, 9, -18, -21, -4, -5, -9, -32, -11, 13, 35, 24, -1, 2, -36, -34, 19, 9, -23, 2, 33, -1, -6, 0, -24, -1, 21, 7},
    '{2, -1, -37, 11, 13, 26, -11, 9, 48, 6, 10, 22, 35, 23, 18, -3, 13, -25, -22, -8, -13, 3, 6, 1, 1, -1, -24, -33, -1, 13, -2, -12, -8, -23, 30, 23, -3, 2, 3, 11, 3, -7, -9, -3, 12, 13, 27, 15, -46, 13, 25, -9, -19, -16, -4, -6, 7, 3, 13, 14, 17, 4, 0, -13, -38, -9, 11, -2, -22, -21, -1, 0, -7, -11, -3, 0, -3, -27, -48, -13, -17, 2, 5, -2, -18, -19, -4, -1, -9, 0, 4, 5, -12, -38, -32, 8, -17, -10, 2, 4, 5, -3, -5, -6, -11, 1, -2, -6, -22, -18, -13, -23, -17, 6, -5, -3, -1, -4, -8, -6, -15, 0, -2, -7, -11, -5, 11, 8, -26, 38, 8, 1, 8, -1, 5, 6, 5, 11, -1, -20, -14, -18, 35, 80, -4, 25, -2, 15, 23, 18, 13, 9, 22, 26, -6, -3, 12, -11, 30, 93, -9, -1, 16, 22, 11, 10, -8, -11, 14, 9, 6, 10, 1, 9, 29, 57, -10, -10, 1, 14, 10, -3, -16, -20, 12, 26, 26, 15, 4, 9, 17, 57, 15, 2, 10, 15, 3, 0, -11, -22, -12, 6, 19, 17, 17, 23, 20, -5, 20, -21, 0, 14, -6, -4, -7, -23, -29, -11, -2, 13, 20, 13, -6, -7, -5, -51, -46, -21, -20, -23, -26, -40, -33, -21, -21, -22, -4, -10, -30, 25, 0, -1, -9, -10, -31, -52, -40, -36, -14, -18, -49, -47, -21, -32, -51, 9},
    '{-3, -2, 32, 4, 13, 1, 4, -8, -15, 26, -11, -61, -29, 3, 28, -1, 28, 39, 24, 2, 18, 25, 29, 19, 16, 15, -8, 30, 36, 43, 64, 46, 35, 55, 1, 11, 13, 11, 1, -11, 2, 6, -5, 3, 10, 12, 35, 41, 30, 40, 4, -10, -11, -26, -36, -38, -36, -16, -10, -16, 1, -23, -21, 6, 42, 20, -5, -4, 4, -9, -15, -14, -14, -11, -3, -7, 1, -14, -34, -17, 23, 2, 25, 21, 20, 21, 34, 44, 37, 16, 0, 0, 1, 12, 13, 26, 44, 31, 32, 18, 17, 27, 35, 40, 25, 1, 3, -3, -2, 25, 33, 67, 30, 15, 7, -7, -13, -2, -17, -23, -7, -1, 2, -7, -6, 14, 13, 31, 15, -12, -18, -17, -22, -8, -3, -7, -3, -11, 6, 13, 5, 15, -11, -26, 1, -33, -15, -3, 4, 14, 0, 3, -12, -23, -1, 9, -7, 1, -14, -23, 52, 24, -13, -2, 10, 7, 3, -4, -12, -4, 6, 10, 11, 12, -2, 29, 34, 1, -1, -8, 5, 7, 3, 8, -1, 2, 11, 4, -1, 6, -10, 23, -8, -18, -29, -27, -9, 2, -4, 9, 4, 0, 10, -6, -17, 5, -17, 23, 4, 4, -3, -19, -27, -14, -7, 3, -4, 2, -6, -30, -23, 9, 7, -9, 2, 14, 0, -9, -8, -18, 0, 12, 0, 4, -3, 6, -18, -3, 26, -37, 1, -10, -36, -30, 4, 15, 22, 24, 25, 13, 21, 46, 6, 7, 47, -1},
    '{-3, 4, -17, 29, 28, 34, 33, 12, -14, -18, 31, 49, 69, 55, -15, 0, -28, -30, 14, 43, 19, 24, 34, 12, 25, 21, 7, 5, 19, 18, -9, -3, -28, -20, 31, 22, 8, 18, 5, -6, -10, 7, 12, 22, 12, 7, -3, 9, -20, -21, 24, -3, -10, -6, -16, -28, -15, -1, -2, 4, 2, 18, 10, 0, -18, -10, 33, 5, -17, -26, -23, -9, -7, -6, -10, -7, 0, 1, 6, -1, -26, 5, 18, 2, -16, -8, -7, 2, -9, -7, -12, 3, -10, -27, -22, -34, -20, -27, -11, 3, -1, 3, 1, -15, -20, -13, -9, -5, -19, -18, -16, -65, -11, -26, -22, 8, 17, 12, 3, -3, 4, 9, 7, 6, 1, 13, 0, -48, -19, 8, -10, 19, 27, 18, 5, 16, 16, 18, 18, 4, 4, -1, 11, 17, 11, 44, -8, 1, 23, 16, 19, 21, 18, 9, 1, 5, -2, 2, 33, 21, -42, 11, 1, -5, 11, 7, 5, 14, 14, 1, -4, 0, -3, 12, 12, -17, -55, -18, -6, -19, -4, 4, 5, -2, 13, 13, 8, 0, 8, 10, 1, 28, -5, -4, -3, -24, -16, -3, 0, 7, 13, 7, 6, 7, 14, -1, -11, 30, 11, -4, 2, -2, -4, 0, -6, 1, 2, -12, 4, 18, 20, -3, -17, 9, 13, -11, -34, -30, -15, -2, -20, -17, -4, -20, -17, -11, -14, -13, -39, 28, 3, 20, 5, 6, -2, -21, -1, -8, -3, -14, -16, -27, -31, -25, -57, 4},
    '{4, 0, -4, 0, -6, -6, -21, -25, -13, 3, 21, -1, -15, 9, 22, -3, 24, 31, -13, -41, -53, -29, -20, -19, -52, -30, 16, -7, 18, 47, 23, -8, 25, 13, -17, -24, -32, -18, 8, 18, 7, 17, 25, 18, 28, 33, 44, 28, -11, -20, -17, -13, -10, 3, 11, 6, -3, 0, 9, 15, 17, 10, 26, 12, -8, -15, -13, -6, 9, 8, -8, -13, -12, -8, 1, -6, -3, 7, 4, 11, 29, 5, 9, 22, 13, 10, 13, 12, -11, -18, -2, -3, -17, 2, 2, 19, -1, 0, 23, 46, 36, 28, 26, 31, 8, -12, -2, 18, -6, -11, 17, 26, 13, 18, 13, 21, 12, 5, -3, 0, -9, -15, 7, 22, 5, -3, 11, 44, 17, 14, -12, -31, -44, -42, -17, 9, -2, -10, -3, -7, -5, 7, -6, 43, -17, -2, -56, -58, -39, -7, 19, 25, 5, -8, -2, -3, 0, 14, -2, 17, -1, -38, -30, -11, -1, 17, 25, 4, -15, -12, -19, -10, -2, 3, 2, -14, -1, -37, -28, 8, 21, 19, 14, -9, -7, -7, -12, -7, -13, 3, 7, 6, 2, 12, -5, 11, 13, 13, 4, -3, 3, 1, -7, -8, -16, 4, 7, -13, 16, 22, 8, -1, 0, 8, 16, 17, 2, 3, 3, 9, -9, 17, -4, -41, -13, -14, -57, -14, -15, -2, 16, 11, 8, 16, 28, 37, -7, 9, 27, -27, 1, -4, -42, -24, -2, -17, 13, 6, 3, -13, -15, 5, -23, -10, 27, 7},
    '{1, -2, 18, -24, -38, -11, 15, 1, 13, -5, -35, -29, 3, -5, -1, -1, -7, 5, -4, -28, -34, -11, -22, -14, 8, 8, 1, 6, 13, 18, 9, 2, -12, -27, -18, -12, -10, -26, -18, 0, 2, -3, -4, -5, 1, 11, -1, 1, 16, 19, -4, -5, -13, -18, 2, 13, 1, -4, 7, 4, 9, -7, -31, -63, -7, 35, -16, -6, -3, -7, 2, 8, 1, 9, 13, 8, 17, 9, 1, -47, 33, 33, -5, 13, 4, 7, 2, 3, 22, 1, 8, 7, 8, 9, -4, -27, 51, 29, -1, 20, 18, 14, -5, 2, 1, -10, 0, 6, 13, 22, 1, -23, 48, 27, 18, 21, 28, 16, -16, -23, -22, -6, 9, 11, 14, 13, 0, -31, -19, 4, 1, 10, 17, 11, -2, -16, -15, -4, 13, 19, 13, -1, -7, -34, -31, -27, -4, 10, 18, 10, 12, -7, -9, 0, 2, -7, -5, -13, -24, -20, 27, -37, -14, -2, 16, 13, 6, 3, 0, -3, -1, -10, 0, -8, -36, -3, 31, -13, -1, -3, 5, 4, 3, 12, -4, -10, -2, 2, 0, -7, -12, -19, 19, 1, 12, 5, 5, 0, 8, 7, -5, -4, 1, -2, -8, -11, -5, -41, -21, -12, -2, 3, 0, -8, -8, -8, -14, 1, 3, -3, 8, 7, 5, -34, 21, 3, 29, 19, 10, 11, 17, -2, -6, 4, 5, 27, 21, 5, -11, -13, 0, 34, 58, 65, 58, 33, 15, 51, 57, 33, 27, 33, 64, 35, 0, -3},
    '{-4, -2, -1, 24, 26, 0, 4, -37, -47, -2, 15, -6, 31, 25, 8, -2, -25, -21, 34, 29, 9, -15, -36, -30, -30, -7, 13, 18, 32, 31, 5, 13, -24, -12, -1, -5, -5, -15, -2, -9, -7, 9, 15, 11, 12, 21, 32, 36, 1, 0, -23, -34, -10, 4, 7, 2, 9, 16, 20, 27, 11, -6, 29, 29, -27, 4, -24, -17, -1, 4, -1, 0, 8, 17, 17, 11, 9, -5, 14, 16, -30, -15, -8, 1, 2, 6, 6, -3, -7, -20, -27, -16, -10, 2, 14, 5, -36, -6, 21, 23, 13, 12, 2, -1, -1, -23, -27, -19, -12, 25, 49, 30, -19, 16, 14, 4, -11, 9, 6, 11, 10, -9, -6, -4, 2, 17, 18, 31, -33, -31, -19, -2, -16, -4, 16, 19, 11, -3, 0, -5, -15, -17, -21, -17, -35, -7, -9, 0, -6, 11, 24, 11, -7, 3, -3, -16, -25, -19, -12, -14, -13, -30, -9, 9, 5, 18, 29, 13, -12, -2, -11, 2, -14, -25, -26, -29, -7, -49, -27, -3, -2, 15, 8, 5, -7, -17, -10, 5, -13, 6, 15, -3, -4, -1, 10, 2, 4, 15, 9, 5, 3, -7, 0, -3, -12, 6, 24, 5, 6, 40, 30, -6, -2, -5, 1, -2, -7, 0, -14, -13, -12, 14, 34, 7, 0, -1, -49, -8, 2, 0, 21, 24, 15, 20, 16, 25, -8, -1, 19, -34, 1, 31, -9, 0, 27, 14, 38, 52, 47, 36, 32, 26, -7, 3, 49, 7},
    '{-3, 0, 21, -16, -20, -22, 7, 19, -8, -14, -9, -11, -26, -18, -26, -1, -2, 20, 48, 25, 11, -9, 2, 22, 23, 6, -4, 18, -8, -29, -20, -24, -33, 3, -15, -22, -16, 8, 16, 9, 8, 2, 7, 11, 1, -20, -22, -34, -2, -54, -43, -26, -14, 2, 11, 10, 1, -10, -5, -2, -6, -13, 2, 12, 1, -59, -51, -18, -12, 5, 18, 6, 11, 8, -2, 0, -3, -18, 28, -6, -15, -49, -32, -8, 9, 15, 23, -11, -12, -6, -17, -15, -8, -15, 52, 17, -19, -52, -29, -5, 13, 18, 12, -6, -6, 20, 23, 1, -11, -4, 21, 28, -13, -40, -6, 11, 16, 9, -3, -17, -14, 6, 19, 14, 0, 15, -4, -3, -16, -42, 11, 17, 23, 10, 3, -20, -25, -1, 8, 9, 14, 16, 18, -18, -33, -14, 12, 6, 4, -2, -5, -32, -26, -10, 2, 9, 3, 15, 9, -32, -8, 21, 17, 18, 10, 6, -6, -25, -4, 0, 12, 19, 6, 9, 11, -52, -6, 5, 23, 18, 14, 20, 10, 1, 2, 6, 13, 11, 6, 11, 25, -24, -47, -42, 10, -6, -7, 0, -4, 8, 12, 15, 14, 8, 17, 0, 12, 14, -26, 4, 20, -11, -36, -23, -3, 9, 22, 16, 9, 2, 4, -3, 10, 22, 6, 19, -2, -11, -19, 0, 5, 25, 9, -4, -2, -5, 17, 20, -2, -22, 3, 18, -2, -11, -20, 10, 11, 4, 4, 9, -26, -17, 36, 36, 11, -13},
    '{-3, 2, 3, 10, 30, 16, 6, 22, 36, 42, 41, 24, 7, 11, 21, -3, 22, 23, 3, -19, -2, 32, 11, 29, -3, -1, 15, 1, -15, -8, 17, 11, 22, 38, -1, -10, -9, 8, 21, 5, 10, 7, 18, 10, -6, -9, 0, 16, -28, -20, -31, -14, 3, 11, 35, 23, 32, 15, 10, -9, 4, -10, -7, 20, -19, -21, -24, -5, 15, 21, 22, 26, 28, 0, -12, -19, -14, -12, -32, 14, -29, 0, -17, 4, 11, 14, 11, 5, -13, -18, -7, -15, -26, -15, -18, 0, -45, 12, 2, 11, 7, 1, -19, -19, -15, -16, 10, 6, 0, -6, 4, 1, -60, 26, -19, -7, 6, 1, -20, -10, -5, -18, 13, 6, -1, -11, -9, -11, -40, -21, -46, -20, 0, -7, -8, 3, 0, -19, -11, -15, -3, -4, 17, 4, -18, -8, -23, -21, -7, -3, -1, 15, -3, -14, -26, -13, 9, 21, 17, -20, 16, 15, -16, -20, -10, -1, 1, -4, -19, -13, -18, 2, 11, 15, -16, -29, 21, 6, -12, -14, -3, -6, -19, -13, -5, 13, 22, 37, 38, 34, 4, 41, 4, 21, 23, 1, 11, 4, 3, 14, 26, 33, 29, 29, 25, 20, 4, 19, -8, 27, 26, 20, 26, 6, 20, 26, 22, 28, 23, 16, 10, 22, 13, -17, -18, -12, -38, 8, 24, 21, 20, 28, 18, 13, -1, 8, -20, 2, 45, -17, 2, -23, -53, 1, -18, -29, 14, 7, -15, -4, -11, -27, -45, 6, 46, 2},
    '{1, 5, 5, -10, 12, 2, -20, 7, 84, 115, 86, 47, 16, 22, -3, 1, 23, 22, 41, 31, 12, 4, -1, -4, -1, 10, 11, 27, 7, 14, 26, 24, 35, 51, 26, 9, -9, -1, 20, -7, -3, 0, 7, 9, 4, 1, -15, 19, 44, 44, 20, 7, -15, -5, 10, 7, 2, 6, 6, 2, -6, 2, 22, 39, 22, 39, 17, 4, -3, -22, 0, 5, 13, 6, -12, -6, 1, 13, 18, 38, -23, 19, -18, -19, -7, -29, -21, -4, 10, -7, -29, -31, -21, 2, 25, 5, -27, 23, -16, -18, -10, -16, 4, 16, 6, -12, -7, -18, -45, -52, -37, 6, -19, 19, 13, 28, 14, 19, 9, 12, -4, -14, -4, 4, 6, -12, -28, -10, 28, 1, 5, 6, 1, 11, -6, -10, -8, -9, -4, 13, 21, 2, -4, 13, 27, 14, -1, -19, -39, -33, -18, -7, -14, -3, 17, 14, 10, -11, 0, 24, 21, 38, 7, 12, -3, -17, -19, -17, 3, 14, 10, -7, -8, -22, -9, 6, -4, 8, -1, 21, 15, 13, 26, 37, 36, 22, 7, -9, 9, 29, 31, 32, -25, -31, -18, 0, 22, 29, 24, 20, 19, 8, 0, 1, 13, 34, 10, 34, 16, 3, -3, -6, 2, 23, 19, 3, 9, 3, -6, -4, -12, -10, -7, 34, -26, 7, 26, 13, -1, -10, -33, -14, -2, -14, 4, -43, -28, -24, 14, 21, -1, 8, 21, 11, -26, -42, -23, -7, 6, 1, -34, -39, -22, -10, 6, 4},
    '{0, -1, 29, -1, -6, -14, -3, -27, -32, 6, -9, -16, -1, 17, 12, 0, -24, 23, 27, 18, 51, 32, 46, 14, 13, 16, 4, 17, 13, 6, 36, 50, -18, 6, -10, -2, 4, -4, 6, -11, -3, -6, -3, 10, -4, -16, -16, 29, 38, 21, 1, -13, -4, -2, -11, -8, -5, 6, -4, -2, -4, -4, 4, 28, 60, 27, -11, -24, -4, -1, 2, -3, 0, 9, 2, 6, -5, -2, -1, -1, 34, 9, 8, -10, 1, 2, -8, -17, -3, 5, 12, 4, 1, 13, 7, 13, 16, 12, 18, 8, 6, 3, -22, -16, 11, 6, 15, -6, -4, 11, 10, 33, 6, 3, 2, -2, -11, -1, -11, 8, 25, 6, 2, 0, -16, -9, 5, 41, -5, -32, 6, 13, -5, 4, 10, 14, 2, -5, 6, 21, 2, -8, -7, 0, -4, -11, 27, 15, -4, -13, -5, -3, -18, -4, 24, 14, -16, -27, -29, -2, 27, 8, -8, 7, 10, 3, 16, 9, -3, 13, 10, -17, -24, -34, -30, 36, -1, -14, -7, -6, -1, 7, 13, 17, 11, 9, 2, -23, -29, -36, -19, 17, -15, -15, -20, -21, -12, -6, -2, 15, 11, 9, -15, -27, -45, -43, -6, 26, 28, 37, 16, -9, 0, -3, -2, -6, -7, -23, -43, -53, -54, -20, 13, -17, -1, 34, 35, 9, 11, -9, 5, 7, -11, -10, -34, -23, -19, -18, 8, -5, 3, 8, -27, -22, 1, 22, 37, 30, 26, 26, 25, 39, 24, -4, 27, 5},
    '{-3, 3, -3, -10, -14, -49, -50, -60, -44, -5, 20, 13, -13, -8, -6, 0, 3, -7, -12, -13, -42, -57, -61, -42, -33, -31, -29, -38, -24, -30, -14, -3, 21, 28, -2, -5, -23, -25, 4, 0, -9, -6, -5, -14, -5, -2, 8, 1, 12, 10, 12, 18, -2, -1, 13, 4, -2, 5, -2, -15, -10, -2, 1, 7, -2, 10, 2, 17, 3, 4, -9, -2, 7, 8, -6, 0, 3, 0, 17, 6, -12, 8, -8, 10, 18, 18, -6, -18, -18, -2, -7, -10, 10, 6, 31, 17, -38, -22, -11, 2, 13, 18, 6, -3, -6, 0, 7, -4, 1, -4, 14, 28, -23, -44, -12, 25, 27, 20, 42, 31, 12, -12, -2, 0, 1, 1, -24, -31, -6, -60, -31, 2, 14, 28, 33, 32, 10, 0, -7, -14, 10, 14, -1, -22, 18, -11, -72, -67, -56, -39, -8, 14, 4, 2, -2, -2, 13, 26, 7, -47, -14, 27, -28, -25, -37, -56, -55, -44, -19, 2, -5, 1, 0, -5, -16, -73, -21, 28, 14, 19, 12, 21, 14, -1, -11, -1, -2, -2, 7, 1, -12, -40, -10, 4, 18, 9, 12, 10, 10, 7, 1, -4, -7, 1, 11, -11, -40, -33, -19, 32, 41, -10, 7, 10, 12, -6, 3, -5, -2, 6, 4, -19, -37, -36, -18, 10, 8, -7, 4, 9, 6, 8, -1, -2, -11, -12, 9, 15, -3, -29, -4, 22, 37, -2, -22, -5, -9, 7, 13, 9, 3, -31, 1, 13, 40, -6},
    '{-1, -2, -39, -18, -18, -8, -9, 9, 14, -44, -39, -21, -8, -27, -1, 2, -6, -38, -16, -25, -20, -27, -11, 1, -11, -33, -4, 17, 5, -33, -20, 28, -13, -6, 0, 14, 6, -6, 7, 17, 5, -5, -9, 2, 2, 18, 30, 15, -4, 10, 12, 6, -7, 7, 5, 1, -6, -10, -8, -16, -19, 1, -4, -31, -2, 21, 1, 11, -5, 4, -2, -8, 8, 0, 1, -7, 0, 14, 14, -3, 2, -4, -12, -2, -3, 9, -13, -24, -12, 6, 16, 11, 1, 7, 47, -8, -19, -17, -7, 14, 16, 23, 7, -30, -44, -18, 12, 4, -9, 5, 15, -14, 3, 4, -6, 13, 15, 20, 18, -15, -40, -26, 14, 7, 10, 0, 5, -11, -5, 8, -2, 10, 18, 27, 31, -10, -50, -20, 21, 11, -1, -15, -13, 19, -8, 0, -6, 1, 4, 17, 13, -24, -42, 8, 18, 3, -3, -26, -16, 15, -5, -17, 14, 21, 7, -13, -31, -23, 3, 17, 21, 0, -10, -13, 5, 25, 31, 17, 8, 17, 10, -22, -25, 1, 3, 13, 25, 4, 4, 1, -3, -7, 28, 22, 13, 2, -13, -12, 1, 10, 3, 8, 10, 3, 17, 21, 21, -30, 22, 30, 17, 13, 4, -2, -5, 1, 2, 3, -7, -4, 12, 23, 23, -13, 28, -3, -23, -13, 0, 6, -13, -8, 12, 19, 19, 5, 17, 25, 2, 32, -1, -5, -2, -6, 13, -3, 10, 29, 12, 0, -23, -32, -17, 1, -31, 7},
    '{1, 4, -7, 6, 5, 2, -8, -2, 11, 40, 19, 11, 24, 20, 13, -3, 30, 34, -30, -23, 6, 15, 19, 15, -7, -14, -7, -21, 12, 35, 14, 2, 42, 29, -8, 0, 7, -10, 9, 11, -4, 2, -6, -4, 9, 9, 10, 17, 1, -2, 1, 2, -12, -12, 2, 0, 2, 2, 3, 4, -3, -4, 10, 4, 26, -12, 0, -10, -12, -3, -4, 0, 4, 7, 6, 5, 2, 9, -1, 9, -8, 11, -13, -16, -1, 4, -6, 1, 13, 19, 6, 3, 14, 26, -11, 6, -23, 20, 20, 1, 7, -4, -12, 1, 24, 0, -4, 2, 5, 16, 4, 21, -33, 19, 0, 5, -2, -6, -18, 11, 15, -9, -1, 2, -2, -24, -12, 31, -28, 4, -17, -6, -4, -3, -2, 24, 14, -2, -5, -21, -29, -47, -34, 10, 12, 14, 5, 3, 8, 1, 1, 19, 6, -5, -10, -23, -23, -12, -3, 2, -33, -3, 8, 7, 3, 5, 3, 6, -8, 5, -4, 0, -4, 7, 5, 6, -30, -5, 1, 7, 4, 10, -15, -13, 2, -2, 4, 15, 13, 21, -1, 20, 39, 54, 9, 24, 19, 2, -6, -8, 3, -2, 9, 17, 9, 9, -1, 14, 31, 44, 24, 12, 17, -1, -1, 1, -1, 4, 2, 4, 7, 13, 9, -5, 1, 14, -38, -12, -10, -5, -1, 2, 5, 9, -6, -14, -33, -26, 15, -17, -2, -9, -51, -39, -2, 3, 10, -4, -8, 8, 12, -16, -49, -38, 36, 3},
    '{3, 0, 20, -14, -18, 8, 12, -25, -52, -35, -19, -9, 44, 18, 3, 2, -25, 7, -12, -4, 43, 25, 48, 25, 17, 4, -4, 0, -3, -1, -13, -13, -24, -4, 10, -1, 9, -1, 7, 2, 2, 6, -3, 2, -17, -34, -25, 32, 23, 16, 14, 15, 10, -2, -9, -6, 1, 8, -2, -6, -19, -3, -3, -5, 39, 44, 40, 9, 10, 2, -14, -3, 4, 7, 16, 3, -15, -14, -9, 5, 25, 53, 24, 0, -1, -11, -26, -13, 2, 20, 16, 15, 2, -12, -39, 23, 7, 42, 6, -3, 0, -7, -12, -4, 5, 0, -4, -8, -17, -12, -33, -4, -8, 19, 7, 2, -10, 8, 8, 19, 20, 1, -2, 2, 7, -16, -19, 12, 7, 16, 16, 6, 4, 14, -2, 12, 19, -6, 13, 30, 29, 1, -2, 12, 25, 13, 35, 15, 42, 19, 1, 27, 6, -6, 9, 19, 18, 13, 8, 19, 13, 16, 2, -16, 6, 1, 7, 26, -7, 5, 12, 13, 15, -7, -48, 9, -29, -9, -5, -19, -20, -10, -22, -9, -5, 3, 0, 8, 10, -49, -88, -20, 0, 13, -14, -8, -13, -21, -5, -1, 5, 9, -6, -5, -10, -51, -84, 5, 24, 22, 9, 9, 1, -13, -9, -6, 0, -5, -10, -15, -20, -34, -53, -8, 17, 27, 43, 19, 10, 7, 6, -6, 2, -9, -20, -25, -16, -28, -41, -26, -3, 2, -15, 3, 24, 48, 33, 11, -6, 17, 37, 2, 13, -26, -10, -8},
    '{1, 3, 33, 27, 31, 28, 36, 1, -8, 7, 49, 51, 46, 44, -12, -3, -29, 5, 40, 47, 17, 34, 43, 20, 17, 6, -29, -24, 0, 55, 29, 24, -27, -31, 24, 18, 20, 30, 11, -3, -6, 16, -13, -19, -22, 24, 30, 44, -30, -30, 23, 1, 11, -11, -6, -13, -22, -26, -26, -6, -9, 12, 23, 23, 16, -24, 12, 3, 9, 5, -4, -17, -23, -26, -10, 6, 11, -6, 9, 17, 3, 10, 3, -5, 17, 19, 4, -21, -22, 13, 11, 22, 7, -12, -10, -28, -4, -4, 2, -12, 5, 14, 6, -18, -20, -3, -3, 5, -12, 4, 26, -53, -31, -2, 0, -3, 2, 12, 6, 4, -10, -5, 13, 10, 11, 22, 21, -35, 2, 13, -2, 9, 14, -7, -11, 19, 23, 8, 11, 5, 2, 9, 24, 0, 20, 33, -15, -9, -13, -30, -7, 29, 25, 2, -2, -1, 1, 9, 36, -8, -45, 20, 8, -18, -29, -28, 19, 36, 13, 6, 9, -8, -14, -2, 17, -23, -34, -10, -35, -28, -20, -10, 30, 23, 10, 4, 6, -18, -8, -12, -9, 15, 8, 1, -34, -24, -4, 5, 11, 14, 8, 7, 14, 9, 14, -7, -3, 49, 1, 1, 3, -45, -44, -31, -25, 5, 2, 8, 2, 3, 0, -12, -23, 41, -20, -24, -8, -39, -51, -29, -22, -21, -14, -15, -11, -25, -11, -8, -41, -16, -2, -23, 0, -2, -24, -59, -33, -56, -100, -68, -23, -55, -59, -21, -26, 7},
    '{0, -3, -10, 8, 6, 8, 8, -31, -26, 1, -14, -48, -26, -14, 12, -2, 27, 15, 10, -4, -25, -22, 2, -31, -59, -56, -46, -71, -47, -4, -16, -31, 31, 13, -20, -6, 16, 15, 23, 20, -7, -37, -36, -32, 2, -4, 20, 30, -16, -4, -14, 2, 13, 20, 11, 13, 12, 7, -13, -27, -9, -11, 33, 18, -49, 13, -11, -22, -11, -3, -14, 12, 26, 10, -13, -22, -17, -5, 28, 29, -20, 7, -11, -10, -10, 0, 5, 8, 17, 2, 5, -23, -34, -7, 18, 52, -14, -8, -14, 16, 3, 11, -1, -19, -2, 25, 26, 0, -26, -23, 6, 18, 0, 0, -26, 1, 4, -4, -26, -10, 26, 33, 34, 4, -21, -26, -9, 5, -38, -18, -44, -9, -5, -16, -11, 11, 17, 20, 12, -22, -22, -9, -13, -3, 22, 4, -12, -21, -13, -4, 8, 2, -5, 6, -23, -38, -24, -8, 6, 0, 31, 15, -7, -14, -2, 6, 16, 9, -9, -10, -23, -15, -12, -4, -5, 42, -12, -28, -13, -15, -7, 1, 7, 6, 1, -1, -13, 2, 2, 11, 1, 35, 0, -24, -13, -26, -8, 14, 12, 9, 13, -4, -17, -3, 6, -1, -9, -4, -22, -30, -22, -12, 2, 5, 7, 6, 1, -5, 1, 16, 22, 14, -3, -25, 23, -33, -3, 15, 10, -11, -8, -16, 2, 1, -1, 1, -15, -11, -2, 3, -2, 9, 30, 36, 29, 31, 31, 13, 21, 4, 17, -5, 2, -14, -18, 7},
    '{-3, 0, -8, -14, 7, 31, 20, 4, 6, -18, -76, -64, -29, 4, 10, -2, 32, 13, -8, 4, 24, 30, 39, 35, 4, -14, -30, -39, -46, 14, 9, 4, 32, 39, 34, 17, -10, -11, 9, 13, 12, 12, -3, -18, -24, -30, 9, 6, 31, 11, 9, 4, -13, -6, 6, 9, 5, 1, -4, -23, -32, -53, -8, -5, 20, 10, 30, 10, 7, 18, 1, -2, 7, 9, 7, -17, -47, -57, -30, -9, 0, 3, 36, 2, -10, -32, -46, -17, 29, 44, -1, -31, -46, -29, -34, -5, -2, 12, -18, -46, -49, -45, -4, 18, 37, 5, -33, -33, -27, -29, -13, 20, -10, 13, -29, -22, -9, 16, 19, 14, 11, -11, -17, -10, -5, -14, 21, 17, 16, 29, 4, 6, 9, 17, 10, 6, 4, -2, -5, 8, 17, 22, 12, 21, 22, 1, -2, 3, 20, 9, -4, 2, -2, 4, -11, -5, 15, 26, -3, 25, -6, -15, -8, -7, -4, -9, -18, -5, -6, -5, -6, -7, 24, 19, 3, 40, -33, -13, -18, -7, -3, -1, -11, 7, 8, -12, -4, 0, 1, 3, 6, 51, -12, 31, 3, 4, 4, -2, -1, 4, 1, -4, -12, -8, -12, 1, 4, 6, 8, 38, 38, 10, 2, -1, 8, 5, 4, -13, -14, -20, -24, -8, 5, 17, 24, 20, 36, 22, 24, 24, 23, 17, 16, -6, -12, -33, -17, 19, 17, 24, -3, -12, 8, 3, 20, 21, 22, 22, 37, 17, 14, 13, 4, 9, 11, 0},
    '{3, -2, 33, -11, -1, 26, 44, 29, 6, 2, -1, 54, 42, 20, 7, 2, -5, 24, 27, 23, -5, -5, 2, 44, 39, 13, 6, 1, -5, 20, 10, -2, 1, 5, -1, 1, -7, -8, -1, 6, 7, 2, 7, -10, -18, -20, -33, -31, 37, 17, -7, -2, 1, -8, 5, 17, 13, -4, -9, -19, -15, -53, -62, -34, 28, 13, -10, 6, 13, 10, 18, 12, 4, -11, -1, -3, -4, -36, -32, -41, 32, 0, 26, 28, 21, 21, 16, -18, -3, 1, 12, -1, 4, -15, -4, -38, 54, 23, 14, 19, 12, 9, -2, -21, 0, 34, 28, 12, 14, 6, -9, -8, 43, 13, 17, 18, 10, 5, -11, -33, -7, 24, 9, 0, 7, 0, -26, -47, 34, 10, 11, 9, 8, -1, -7, -23, -12, -4, -2, 19, 15, 3, -21, -38, -20, -23, 11, 12, 1, -11, -16, -29, -13, -2, 1, 2, 1, -14, -32, -14, 32, -1, -8, -10, -11, -4, -9, -25, -2, 1, 9, 3, 2, -18, -16, 7, 14, -15, 1, -13, -18, -23, 9, 10, -3, -7, 4, -6, -17, -22, -3, -1, -31, -40, -1, -17, -21, -9, 10, 17, 7, 6, -10, -20, -25, -20, 1, -5, -3, -23, -16, -11, -16, -3, 5, -2, -2, 4, -4, -17, -21, -15, 0, -23, 19, 21, -5, -34, -10, 4, -8, -10, -9, 3, -4, 5, 0, -6, 5, -5, -2, 14, -21, -28, 8, 44, 5, 9, 31, 29, 21, 49, 43, 23, 15, -1},
    '{3, 0, 30, -11, -5, 38, 18, 8, -21, -52, -55, 58, 59, 33, 14, 3, -1, 28, -4, 0, -9, 12, -21, -18, 4, 11, -10, 0, 17, 24, 13, -22, 22, 10, 5, 11, 6, 5, -18, -17, 12, 24, 18, 7, -2, -16, -50, -52, -21, 3, 29, 18, -18, -20, -9, -2, -1, 2, 10, 11, 12, -3, -44, -83, 5, 8, 20, 0, -19, -16, -2, 4, 1, 9, 8, 11, 11, 8, -8, -74, 10, 18, 11, -2, 0, 2, -11, -12, -2, 3, 18, 24, 17, 17, 10, -49, 16, -6, -9, 5, 8, 6, 1, -3, -18, -26, -6, 16, 34, 34, 5, -34, 18, -14, 5, 26, 12, 13, -4, 2, -15, -53, -35, 1, 26, 25, 7, -40, -1, -4, 15, 14, 6, -13, -23, 8, -5, -49, -20, 4, 19, 17, 12, 10, -5, -25, 2, 9, 2, -26, -28, 0, -39, -35, 5, 15, 5, 2, 8, 19, -19, -36, -29, -15, 4, 13, -10, -21, -29, 0, 23, 15, 19, 10, 2, 45, -13, -16, -12, -2, 10, 21, 25, 4, 1, 8, 10, 9, 10, -4, -3, 50, -10, 13, 13, 8, -2, 21, 18, 17, 14, 5, -2, -11, -2, -1, -4, 37, 19, -2, -4, 14, 9, 18, 14, 14, 18, 23, 4, -12, 7, 9, -10, 13, 14, 23, 25, -9, -10, 8, -11, -26, 1, 2, -28, -7, 20, 23, 15, 10, 3, 2, 11, -4, 6, 0, -24, 0, 9, 2, -7, 34, 52, 51, 2, -1},
    '{-2, -3, -3, -10, -22, 0, -25, -47, -66, -51, -37, -27, -14, -10, 5, 1, 27, 19, -10, -21, 0, -2, 6, -19, -38, -57, -56, -20, -10, -18, 0, -3, 30, 43, -3, -11, 7, -5, 10, -6, -12, -22, -30, -27, -44, -40, -3, 6, 2, 29, 0, 4, 1, 0, 0, 8, 14, 9, -9, -32, -52, -64, -34, 6, -32, 27, 18, -13, -16, -7, 1, 24, 29, 23, 3, -18, -35, -70, -53, -13, -31, 18, -1, -3, -5, 2, 7, 6, 21, 19, 17, -1, -20, -44, -44, 5, -9, 32, 11, 21, 5, 2, -7, -16, 5, 4, 10, 5, -2, 0, 11, 25, 3, 17, 5, 8, 8, 3, -11, 8, 16, -2, -2, 0, -3, -18, -28, -3, -5, 12, -23, -9, -3, -15, -19, -6, 1, 6, 0, 3, -1, -11, -33, -6, 21, 15, -3, -9, -8, -15, -20, -12, -4, 10, 13, 0, -10, 1, -12, 0, 23, 18, 9, 9, 4, -7, -11, -7, 5, 15, 17, 6, -2, -7, -8, 35, -32, 0, 5, 9, 6, 6, -9, -12, -13, 0, 10, 14, -6, 9, 10, 9, -6, 19, -4, -2, 0, -1, 6, 2, -4, 5, 3, 2, -8, 9, 5, -37, 11, 27, -13, -26, -20, -18, -2, -5, 2, 1, 5, 3, 3, 23, 14, -36, 23, 6, 15, 6, 8, 3, 1, -1, 5, 10, -2, 16, 5, 6, -10, -20, -2, -2, -5, 11, 28, 47, 42, 51, 54, 35, 36, 25, 33, 6, 5, -6},
    '{-1, 3, 2, -1, -1, 1, 1, 4, 2, 0, -2, -3, -2, 3, -4, 3, 3, 1, -3, -4, -3, 1, 3, 5, -2, -4, 3, -1, 0, -1, -2, 0, -3, -3, -3, 0, 1, -6, 2, -2, 2, 0, 1, -4, -6, -3, -4, -2, 0, -2, 0, -1, -5, -6, -2, 2, -4, -4, 3, 3, 0, -2, -2, -2, -4, 1, 1, 2, -6, 0, -4, -1, -6, -4, 3, 1, -7, -3, 2, -2, -3, -1, 2, -3, -2, -1, -2, -2, -4, 3, 1, 1, -1, -7, 0, 2, -2, -1, -2, -2, -6, -5, 0, 1, -2, -2, -1, -5, -1, 0, 4, 1, 0, -1, -5, -5, -4, -7, 1, 1, -4, -9, 2, 2, 3, -7, 0, -2, 3, -3, -6, 0, -5, -7, 1, -2, -6, -6, 1, -2, 0, -3, 2, 2, 0, 1, -1, 3, 1, -5, -5, -6, -3, -5, 3, 3, 0, 0, -3, -2, 2, 1, 1, -1, 2, -2, 2, 2, -3, -3, 1, -2, -2, 2, 2, -4, -5, 2, -1, 2, -3, 2, -2, -3, 3, -4, 1, -4, -4, 1, -3, -3, -1, 1, -5, 1, -2, 1, -3, -1, -3, -5, -1, -9, -4, -4, -3, -2, -2, -1, -4, -1, -4, -6, -1, -1, -4, -4, -5, 0, -4, -4, 3, 3, -2, -2, -4, -3, -1, 4, 0, 1, -1, -2, -7, -3, -3, 0, -2, 4, -3, 2, 3, 0, -4, 1, -3, -3, 0, -1, -6, -2, -4, 1, 4, -1},
    '{-3, -4, -37, -8, -13, 7, 6, -12, -15, -27, -23, -15, -4, -11, -4, 2, 2, -40, -39, -43, -58, -51, -19, -36, -62, -46, 19, 38, 29, 8, -27, -26, -4, -42, 12, 15, -15, -16, -5, -10, -24, -27, -19, -22, 1, 28, 28, -19, 32, 30, 26, 18, 3, 4, 9, 11, -6, -11, 0, -10, 10, 25, 9, -14, -21, 29, 16, 8, 6, 11, 6, -3, -7, -5, 17, 16, 23, 42, 25, 13, 0, 0, 17, 22, 14, 7, -7, -7, 2, -16, 12, 17, 25, 18, 48, 34, 19, 4, 17, 10, 16, 17, 15, 7, -7, -15, 2, 23, 18, -4, 7, 28, 36, 27, 3, -1, 26, 9, 7, -14, 10, 2, -7, 13, 14, -10, -5, -9, 55, 37, 12, 2, 5, 6, -2, 5, 23, 5, 2, 11, 10, -1, -28, -28, 15, 18, 14, 2, -9, -8, 8, 3, 10, 2, -9, -14, 4, -4, -26, -19, 27, -7, -14, -32, -23, -21, -7, 0, -1, -18, -25, -18, -14, -17, 11, 31, 31, -44, -50, -41, -25, -15, 4, 12, -3, -28, -34, -24, -21, -28, -6, -11, -11, -84, -32, -13, -4, 6, 15, 15, 2, -24, -22, -15, -8, -13, -4, -39, -19, -54, -11, 5, 16, 23, 25, 10, 11, -18, -42, -18, 8, -7, -19, -1, 26, 7, 28, 1, 3, 9, 19, 4, 22, -5, -31, -17, 18, -3, -43, -16, -4, 12, 9, 2, 20, 27, 2, 22, 32, 13, -2, 5, 32, 39, -28, -5},
    '{-2, 2, -24, -24, -22, -28, -12, 2, 24, -5, -6, 18, -6, -17, -17, 0, 26, 2, -33, 0, 32, -3, 2, 9, 10, 5, 15, 21, 6, 16, -16, -46, 31, 22, 22, 10, 15, 7, -3, 3, 9, -1, -2, 15, 18, 13, 11, 9, 18, 0, 0, 19, 9, -1, 0, 3, -3, 0, -6, 15, 4, 7, 2, -3, -10, 18, 4, 1, 2, 0, -3, 1, 0, 2, 3, 14, 7, -4, -12, 13, -1, 15, 4, 2, 13, -2, -6, 9, 14, 3, 9, 10, 19, 8, 3, 44, 0, 31, 17, -3, 13, -4, 3, 32, 18, -3, 10, 7, 1, -4, -3, 24, 19, 15, 13, 3, 7, -7, 6, 13, 16, 4, -7, -10, -17, -24, -1, -3, 45, -11, -4, -13, -5, -4, 2, 13, 17, -1, -1, 4, -4, -11, -14, -21, 17, -7, 14, 0, -5, -11, -24, 3, 9, -14, 14, 5, -4, 5, -25, -32, 9, 27, 2, -5, -6, -16, -13, -3, 5, 7, 10, 8, -8, -13, -12, 5, -37, -5, -5, -6, -8, -2, -8, -1, 7, 4, 2, 3, -17, -32, -16, -4, -15, -14, -21, -3, 4, -13, -1, 1, -4, -5, -3, 5, -18, -49, -42, -32, -5, -18, -1, 5, -6, -17, 0, 3, 12, 14, 8, 5, -34, -48, -38, 11, 25, 25, 51, 11, 4, 17, 11, -2, -1, -8, -22, -19, -41, -46, -45, -20, -2, -7, -26, -29, 8, 58, 20, -18, 3, 1, 39, 10, -28, -31, -1, -5},
    '{-1, 0, 27, 28, 10, 1, 3, -7, -8, 1, -13, -15, 54, 20, -2, 2, -26, 16, 27, -2, -1, -6, -48, -6, -7, -9, -15, -16, 23, 25, -5, 21, -30, -11, -12, -34, -40, -35, -20, 3, 4, 3, 4, -7, 3, -4, 1, 25, -8, 8, -35, -38, -37, -14, 1, -2, 5, 5, 7, -4, 0, -18, -28, -25, 25, 22, -45, -28, -22, -5, 6, 2, -2, 13, 11, -3, -6, 9, 20, -18, 35, 18, -34, -18, -9, 7, 8, 6, 7, 1, -2, -3, -20, 1, 5, -30, 36, 14, -5, 13, 0, 4, -7, 0, 2, -6, -13, -6, 0, 21, 31, -34, 10, 7, 13, 10, 3, 12, 11, 0, -18, -19, -2, 10, 16, 26, 17, -15, -48, -12, 8, 8, 6, 17, 17, 3, -15, -18, -2, -5, 17, 9, 31, 2, -52, -16, -6, 3, 9, 25, 24, 2, -13, 2, -16, -12, 13, 11, 9, 1, -45, -47, 8, 13, 14, 26, 15, -23, -8, 8, -20, -17, 9, 7, -18, -20, 36, -3, 8, 9, 12, 20, 11, -19, 1, 6, -7, 5, 13, 10, -1, 26, 27, 25, 24, 14, 10, 15, 10, 2, 5, -7, -15, -4, -11, -16, 3, 45, -5, 39, 20, 1, 5, 9, 13, 8, 3, -10, -21, -24, -34, -5, -11, -9, 12, -15, -44, -9, -3, 8, 18, 11, 1, -6, -13, 11, -16, 6, 22, -26, 4, 1, 17, 31, 11, -14, 9, 21, 10, 5, 2, 20, -31, -22, 38, 6},
    '{2, 5, 2, 18, 38, 22, 12, 2, 20, 28, 56, 55, 46, 38, 8, 3, 28, 17, 10, 36, 35, 5, 13, 13, 30, 35, 18, 19, 21, 20, -3, -18, 38, 35, 54, 33, 27, 12, 4, 2, 5, 7, -8, -3, 2, -10, -15, -25, 37, 13, 29, 28, 12, 0, 2, 1, 8, 8, -4, -20, -27, -25, -7, -11, 29, -8, 21, -3, -11, -14, -16, -20, -9, -14, -18, -33, -47, -35, -14, -13, 34, -33, 10, -25, -19, -14, -19, 12, 9, -16, -29, -21, -11, -8, -4, -19, 5, 11, 21, 1, 15, 24, 30, 42, 5, -16, -5, 8, 10, 5, -3, 8, 4, 17, 25, 30, 38, 39, 17, 1, -7, 3, 15, 27, 14, 18, 8, 12, 49, 6, -12, 12, 12, 4, -25, -21, 13, 0, 0, 10, 11, 18, -18, -22, 18, -13, -24, -16, -17, -22, -40, -10, 15, -21, -18, -5, 5, 8, -23, -42, -1, -17, 10, -3, -14, -13, -17, 8, 5, 7, -6, -8, 3, 0, -19, -40, -7, -8, -11, -9, -1, 12, 8, 2, 9, 20, 9, -4, -10, 5, -23, -51, 0, 14, -22, -19, -3, 3, -1, -18, 2, 6, 11, 8, -2, -7, -37, -29, -4, 19, 17, 11, 1, 10, 3, -7, 5, 1, 5, 24, -10, -43, -2, 22, 14, 8, 2, 26, 20, 13, 8, 10, 8, -8, 8, 20, 9, -10, 14, 24, -3, -28, -23, 10, 15, -4, 7, -5, -25, -16, -19, 25, 16, 18, 5, 3},
    '{-4, -2, -12, -8, -10, -35, -33, 17, 18, 33, 16, -13, -11, -31, 6, 3, 32, 17, -44, -33, -20, -44, -58, 2, 32, 20, 19, 5, 0, 16, -14, -27, 32, -1, -49, -17, -20, -25, -20, -5, 8, 10, 11, 18, 10, -6, -3, 3, -11, -30, -31, -13, -13, -10, -9, -13, -5, 8, 17, 26, 3, -1, 8, -7, -9, -9, 3, -1, -2, 6, 5, 7, -16, -13, 24, 31, 2, 1, -1, -2, -17, 13, 5, 7, 12, 8, 10, -10, -39, -8, 37, 38, 21, 11, -26, 20, -8, -6, 4, 1, -1, -11, -18, -28, -3, 30, 35, 30, -1, -20, -36, 4, -29, 7, -6, -22, -17, -12, -11, 4, 19, 22, 23, 13, -13, -43, -21, 22, -8, 14, -3, -18, 0, -4, -6, 16, 28, 22, 9, -17, -15, -32, -25, 18, 42, 32, 14, -7, -2, -5, -5, 26, 23, -8, -23, -26, -11, -1, -5, -3, -17, 21, 11, 0, -1, -8, 1, 16, 1, -17, -16, -14, -9, 22, 1, -2, -36, -3, 3, 4, 11, -3, -10, -11, -1, -4, 3, 3, 0, 13, -20, -12, 28, 47, 1, 14, 18, 6, -6, -20, -13, -9, 4, 14, 1, -6, -24, 0, 42, 6, 2, 11, 9, -7, 1, -1, -8, -12, 2, 4, 6, -5, -23, -4, -16, -5, -11, 2, -11, -5, -5, 5, 7, 0, -3, 0, -17, -25, -32, -5, 1, -20, -33, -14, -1, 5, 5, -11, -1, -22, -11, 2, -8, -32, -43, 4},
    '{2, 0, 24, 19, 18, 24, 33, 2, -15, 20, 14, 23, 48, 25, 24, -2, -21, 20, 36, 8, 16, 67, 54, 36, 8, 19, 15, -1, 18, 28, 9, 23, -14, 14, -10, -19, -9, 25, 11, -14, -15, -1, 9, 0, -10, -10, -11, 27, -8, -13, -5, -16, -1, 6, 4, -11, -5, -3, -8, -1, 4, -6, -2, 11, 22, -11, 3, -1, 7, 9, 0, -1, 8, 9, 3, 0, -3, 7, -1, 8, 5, 17, 3, 14, 15, 10, -11, -1, 7, 11, 3, -3, -18, 9, -5, -22, 1, -4, 18, 14, 4, -13, -20, -23, -3, -7, 5, -1, -1, 16, 27, -22, -26, -1, 16, 18, -2, 1, -8, -1, -12, -13, 11, 13, 12, 13, 9, 7, -68, -31, 3, 16, 6, 4, 13, 6, -4, -12, 2, 1, -5, -5, 22, 12, -36, -11, -6, -8, -11, 11, 30, 14, -15, -10, -11, -8, -13, 9, 33, 8, -32, -36, -12, -8, -7, 9, 26, 7, -8, -2, -10, -3, -10, 12, -9, 2, 28, 1, -4, -1, -2, 13, 10, 10, 13, 4, 6, 13, 14, 12, 6, 37, 52, 53, 24, 8, -2, -2, 1, 9, 15, 3, 7, 4, -3, 11, 13, 43, 24, 70, 8, -12, 0, 11, 0, 18, 11, -1, 5, -1, -1, 15, 5, 1, -21, -3, -37, -6, -6, 6, 3, 24, 11, 2, 5, 10, -6, 11, 18, -11, 2, 2, 21, 23, 1, -25, 9, 10, -9, 0, 7, -8, -24, -14, 47, 2},
    '{4, 3, 11, -10, -5, -18, 3, -7, -10, 26, 55, 26, 4, 5, -16, -1, -14, -8, 41, 35, 64, 33, 29, 21, 14, 32, 45, 23, -6, 8, -8, -2, -6, 28, 0, 7, 33, 19, 9, -13, -10, -1, 4, 8, -1, -1, 3, 33, 1, -8, -2, 9, 19, -4, -13, -13, -11, -13, -7, -1, 2, 10, 17, 44, 16, 4, 4, -6, -4, -7, -3, -4, -5, 0, 0, 11, 10, 18, 18, 35, -23, 17, 4, -17, -4, 3, 1, 2, -10, 10, 11, 16, 15, 32, 28, -3, -39, 28, 12, -3, -3, 0, -13, -6, 3, 6, 23, 6, -3, 5, 3, 2, -25, 7, 1, 1, -11, -10, -6, 10, 18, 4, 5, -12, -15, -9, -13, -12, 18, -17, 18, 7, -5, -7, 4, 19, 13, -6, -22, -12, -12, 5, 27, -38, 12, 22, 18, 3, -12, -19, -4, 9, -5, -17, -6, 9, -3, 21, 19, -61, 1, 25, 4, 14, 9, -17, -5, -8, -21, -5, 9, 23, -6, -36, -64, -83, -8, 3, 7, 13, 4, 8, -4, -1, -2, 13, 31, 29, -10, -66, -84, -78, -24, -17, -15, -10, -2, -16, 10, 11, 5, 8, 21, 8, -41, -85, -69, -43, 8, 38, 20, -2, 0, -5, 11, 11, 15, 11, -4, -31, -64, -55, -30, -27, 0, 36, 2, 13, 19, 26, 15, 31, 0, -1, -26, -43, -37, -27, -26, -25, 0, -12, -12, -15, -8, -16, 9, -15, -44, 4, -4, -19, -31, -18, 2, 5},
    '{2, 0, 12, 1, -12, -33, -52, -47, 8, -17, -26, 21, 7, -8, -4, 2, -21, -25, 34, 23, -52, -60, -50, -49, -25, -16, -5, 8, 2, -20, -1, 31, -21, 28, 42, 9, -42, -47, -40, -13, -4, -19, -26, -21, -7, 25, -3, -10, -25, 30, 61, -1, -5, -26, -27, -7, 4, -15, -12, -12, -15, 9, -8, 22, 3, 13, 33, -14, -10, -30, -26, 12, 3, -2, 8, -8, -5, 11, 5, 12, 20, 3, 29, -12, -18, -64, -42, 17, 34, 22, 25, 10, 11, 26, 41, -8, 1, 6, 28, 2, -34, -54, -31, 29, 28, 7, 9, -1, 13, 29, 39, 21, -15, 7, 4, -45, -24, -10, 1, 21, 16, -4, -11, -33, -52, -53, -44, -24, -3, -19, -5, -5, -10, -10, 0, 13, 16, -2, -17, -18, -34, -82, -48, -30, -32, -20, 32, 18, -16, -34, -12, -4, 13, 3, 1, 0, -17, -14, 20, 8, 32, -28, 11, 19, 15, -4, -6, -3, 20, 11, -8, -21, -31, -3, 29, 38, 24, -66, -24, 14, 17, -3, -5, 4, 13, -5, -9, -36, -45, -13, 23, 35, -28, -56, -17, 12, 9, 9, 5, 3, 7, -10, -16, -39, -28, 2, 25, 9, -38, -40, -4, 4, 8, 19, 5, 5, 4, -22, -46, -23, -6, 5, -5, -15, -9, -31, -16, -31, -13, 5, -2, 9, -3, -8, -33, -36, -13, -8, -4, -2, -3, 25, 44, 17, -27, -12, -19, 2, -7, 13, 9, -4, -19, -15, 11, -4},
    '{-2, 3, -29, -12, -11, -30, -9, -22, -35, 2, -24, -49, -48, -29, -15, -1, 25, -9, -38, -47, -66, -68, -84, -104, -68, -40, -8, -35, -5, 2, -24, -36, 19, -1, -26, -30, -37, -32, -11, -9, -17, -14, -12, -27, -6, -7, 8, 18, -12, 2, -11, -11, -12, 10, 12, 4, 2, 4, 6, -5, 5, -23, 2, 3, -31, 13, -7, -9, 4, 16, 2, 5, 6, 7, 15, 2, 2, -6, 3, 10, -9, 18, -1, 17, 10, 12, 6, 11, 20, 10, 15, 5, 4, 5, -5, 42, 23, 32, 15, 20, 13, 12, 14, 13, 12, 8, 5, 11, 12, 15, 3, 31, 44, 41, 35, 9, 27, 8, 5, -5, 3, 12, 15, 1, 5, -10, 6, 37, 5, 29, 5, -3, 7, 4, -1, 4, 5, 15, 8, -4, 3, -18, -10, 25, -13, -10, 1, -7, -1, -1, 1, 12, 10, 20, -1, -21, -7, -12, -17, 5, 39, -19, -30, -19, -9, -8, -2, 5, -5, -8, -7, -10, -6, -14, -8, 15, 46, -4, -29, -29, -14, -17, -16, -1, -10, -9, -11, 1, -14, -9, -2, -23, 38, 4, -9, -9, -1, -8, -2, -1, -7, 1, 1, -2, -16, -17, -8, -52, -23, -29, -7, 6, 6, -5, 7, 2, -9, -6, 0, 4, -2, 1, -6, -34, 24, -2, 27, 4, 4, 1, 3, -11, -6, -7, -6, 27, 6, -8, -25, -24, -3, 2, 8, 24, 41, 43, 3, 21, 36, 18, 30, 38, 47, 14, -7, -3},
    '{3, 1, -17, 5, -5, -5, 26, 4, -11, -40, -17, -8, 26, 10, -22, 1, -27, -44, 36, 28, 5, -3, -7, -12, 16, 8, 4, 8, 25, 12, -11, 4, -35, -28, -20, -14, -11, -2, 7, 1, 0, 2, 13, 10, 11, 29, 18, 33, 10, -4, -9, -27, -6, 11, 4, 7, 5, 13, 15, 9, 11, 16, 15, 29, -11, 17, -3, 0, 6, 13, 3, -7, 6, 3, 7, 3, 12, 22, 46, 2, 9, 12, -6, 12, 14, 15, -6, -19, -8, -28, -20, 2, -4, -1, 48, -31, 33, 2, 6, 10, 15, 22, -5, 4, 3, -10, -11, 3, 3, 3, 7, -27, 21, 12, 11, 3, 9, 8, 3, 2, -4, -2, 8, 15, 19, 19, -2, -32, -2, -4, 5, 10, 26, 15, 13, -3, -4, -3, 12, 10, 9, 1, -4, -36, -19, -19, -11, 3, 17, 15, 21, 3, -6, 12, 7, 3, -4, 0, 2, -33, -18, -28, 1, 1, 11, 5, 10, 5, 0, -2, 0, -2, -7, 1, -16, -17, 13, -34, -1, -11, -7, -3, -6, -3, -8, -12, -7, -2, 3, -8, -14, -28, 5, -15, 7, -4, -9, 4, 9, 2, 3, 2, -2, -9, 6, -7, -3, 3, -19, 4, 16, 4, 11, 2, 1, 5, 0, 10, -6, 0, 0, -3, 0, 12, 21, 7, -5, 2, 6, 14, 18, 13, 8, 7, 6, 17, 26, 29, -32, -28, -4, 8, 40, 36, 34, 8, 3, 37, 13, 13, 14, 0, 54, 50, -19, -3},
    '{0, 5, 41, 28, 34, 48, 36, 5, -9, 35, 73, 80, 78, 51, -4, -1, -27, 30, 45, 37, 10, 23, 25, 11, 13, 17, 14, 14, 31, 37, 5, 13, -6, 4, -15, -5, -7, 11, 6, 1, -5, -4, -2, 3, -4, -8, -19, 9, 48, 11, -25, -19, -11, -17, 6, 17, 15, 1, -10, -15, -21, -11, -6, 9, 56, -44, -48, -23, -5, -16, 16, 24, 15, -17, -18, -14, -26, -25, 2, -1, 51, -26, -34, -15, -5, -23, -13, -1, 3, -14, -9, -12, -6, -20, -18, -23, 2, -46, -31, -15, -11, -29, -26, 6, 7, -8, -5, -1, 21, 10, -9, -29, -28, -11, -36, -21, -15, -7, 2, 29, 19, -6, -1, 7, 7, 21, 6, -24, -22, 59, -7, 0, 1, 10, 19, 19, -1, -6, 2, -1, -4, 4, 2, -12, -13, 13, 2, 11, 20, 21, 30, 13, 3, 4, 11, 1, 2, -4, 19, 0, -20, -9, 11, 13, 15, 22, 19, -1, 6, 8, 12, 2, 7, 8, 25, 10, 21, 23, 11, -9, -4, 23, 24, 5, 3, -1, -6, 3, 14, 4, -5, 42, 9, 8, 4, -20, -4, 12, 11, 7, -1, -2, -11, 7, 14, -21, -27, 36, 30, -5, -4, -15, -11, 5, 7, -5, -8, -2, -23, -20, -22, -43, -45, -10, -5, -27, -29, -14, -49, -10, -3, -31, -49, -39, -72, -67, -20, -35, -16, 36, 2, -13, -41, -42, -32, 8, -18, -62, -69, -71, -86, -47, -33, -25, -4, 10},
    '{4, 0, -38, -16, -27, -38, -53, -58, -48, -22, -28, -65, -57, -35, 0, -3, -3, -32, -45, -60, -91, -83, -87, -107, -54, -15, 7, -14, -4, -4, -16, -5, -1, 6, -11, -30, -53, -78, -51, -55, -29, -11, -3, -24, 12, 25, 9, 17, 35, 28, -14, 3, 3, 9, 9, 6, -6, -9, -14, -2, -9, -11, -13, -9, 13, 30, -6, -5, 2, 0, 2, 10, 1, 5, -7, -1, -15, -13, 7, 4, -34, -2, -11, -8, -1, 4, 16, 12, 6, 16, 13, 5, 10, 12, 17, 29, -45, 2, 9, 2, 5, 7, -10, -10, -15, -7, -4, 7, 16, 22, 16, 50, -31, -3, 19, 5, 10, 4, -18, -8, -8, -20, -12, 8, 8, -6, 17, 65, -59, -6, 8, 8, 28, 39, 23, 17, 3, -1, 3, 7, 7, -16, -12, 31, -27, -21, -16, 10, 18, 33, 51, 52, 19, -1, 1, -2, 12, 2, -18, 4, 29, -37, -60, -19, -22, -31, -4, 14, 2, -5, -12, -9, -10, -27, -44, -17, 4, -16, -31, -19, -22, -43, -56, -27, -8, 8, 8, -7, 1, -7, -31, -31, 12, 23, 27, 8, 5, -2, -6, -10, -2, 8, 1, -5, 9, 16, 8, -41, -4, 27, 39, 17, 18, 2, 10, -4, -4, -18, -13, -1, 10, 29, 23, 12, 20, 11, 37, 12, 6, 3, 11, 10, -7, -10, -4, 26, 26, 24, -7, -36, 1, 6, 30, 27, 12, 27, 32, 46, 46, 42, 37, 40, 57, 25, 24, -16},
    '{3, 2, 16, -23, -34, -35, -16, 2, 5, 11, -45, -95, -100, -49, 9, 3, 12, 25, -9, -36, -22, -20, -4, 16, -4, -6, 5, 5, -21, -19, 11, -5, 9, 7, -39, -35, -18, -21, 8, 14, 11, 1, -4, -15, -22, -35, -17, -2, -2, 14, -30, -22, -10, 1, 16, 10, 15, 13, 10, 7, 2, -27, -18, -7, -19, 9, -25, -6, 1, 3, -1, -5, 16, 19, 17, 9, 10, 3, -11, 5, -12, 25, -3, 14, 8, 14, 3, 4, 23, 10, 17, 1, -8, 5, -8, -5, 6, 29, 16, 14, 6, 3, -5, -7, 8, -4, 6, 5, 1, 13, 23, 18, 19, 16, 8, -7, -1, -6, -7, -8, 10, -1, 2, 10, 4, 2, 1, 31, -29, -22, -19, -10, -8, -10, 3, 6, -1, -7, -6, -2, 1, -8, -11, 8, -9, -14, 11, 3, 2, 0, 8, -1, -18, -1, -1, -17, -22, 8, -9, -2, 20, -5, -13, 9, 8, 11, 20, 6, -7, 4, 6, 1, -14, 7, -18, -15, 5, -20, -3, 4, -2, 4, 1, 0, -9, -6, 4, 12, -1, 10, 18, -5, 13, 7, 8, 10, 0, -12, -7, -3, -2, 0, 0, 1, -16, -10, 12, -15, -9, 29, 7, -24, -9, -24, -10, -11, -6, -4, -8, -5, -7, 17, 22, -11, 26, 12, -3, -1, 12, 12, 14, 21, 16, 17, 6, 29, 5, 2, 7, -37, -2, 7, 13, 22, 57, 42, 42, 61, 71, 51, 47, 49, 38, 9, 29, -6},
    '{1, -1, -7, 15, 5, 16, -2, -34, 13, 30, 19, -1, -14, 22, 23, 3, 30, 27, -6, 6, 21, 11, -15, -39, -46, -31, -31, -33, -31, 12, 18, 19, 23, 37, 22, 8, 8, -19, -37, -28, -24, -33, -62, -53, -17, -17, 12, 29, 22, 40, 40, 31, 21, 8, -11, 11, 15, 1, -26, -10, -7, -45, -48, 30, 46, 35, 44, 18, 14, 19, 24, 25, 15, 5, -2, -1, -4, -38, -81, 29, 46, 14, 39, 17, 18, 29, 20, 16, 17, 5, -1, -6, -4, -2, -21, 32, 15, -21, 11, 13, 5, -10, -28, -49, -15, 6, 6, -4, 3, 3, -1, 0, 2, -11, -29, -42, -54, -50, -35, -18, 1, 4, 9, -2, 4, -10, 0, -11, 20, -11, -38, -21, -28, -1, 24, 17, 11, 1, 19, 14, 12, 7, -5, 4, 9, -32, -28, 17, 6, 0, -3, 10, 10, 1, 12, 6, 3, 4, 17, 22, 14, 8, 12, -11, -10, -9, 7, 16, 11, 8, 16, 0, -12, 3, 19, 63, -1, 40, 25, -12, -19, -17, 12, 11, 14, 2, -16, -5, -16, -33, -19, 40, 20, 11, 5, -8, -27, -11, 5, 7, 4, -10, -13, -6, -14, -22, -13, 6, 20, -41, -2, 25, -1, -8, -12, -3, 3, 5, -8, -11, -10, -11, -2, -16, 8, -2, 7, 5, -6, -2, -3, 0, 9, 7, -1, -10, -24, -21, 25, 28, 1, -19, -41, -34, 10, 19, 18, -7, 2, -7, 26, 34, -31, -50, -2, 8},
    '{0, -2, 19, -29, -28, -17, -11, -5, -5, -21, -52, -47, -33, -15, -17, 0, 0, 15, -7, -40, -16, -1, -7, -23, -38, -47, -63, -54, -41, -6, 14, 6, -16, 2, 0, 7, 10, 10, 16, 6, 2, -11, -15, -35, -16, -3, -25, -35, -10, 42, 14, 20, 17, 18, 19, 26, 13, 5, 9, 3, 6, -19, -20, -16, -15, 40, -3, 17, 17, 4, 0, 1, 13, 13, 19, 10, 16, -13, -7, -12, -6, 13, -7, 16, 1, -8, -6, -4, 17, 20, 6, 0, 14, -1, -29, -30, 36, 24, -11, -2, 5, -2, 0, 2, -5, -15, -1, 8, 19, 8, -34, -45, 32, 17, -1, -6, 12, 1, -13, -21, -23, -17, 6, 22, 18, -5, -20, -40, -2, -7, -11, -9, -2, -6, -11, -5, -11, -9, 19, 34, 16, 1, 10, 4, 7, -16, -10, -6, -11, -14, -9, -11, -20, -2, 16, 5, -5, 0, -4, 9, 25, 7, -24, -12, -1, -6, 2, -11, -10, 14, 13, -8, -14, -4, 1, 36, 23, -2, -9, -13, -5, 1, 0, 5, -2, 4, -3, 2, -18, -12, -2, 10, 4, 1, -6, -6, 6, 3, -5, 11, 8, 10, -4, -27, -24, -14, -5, -26, -20, 4, 0, 11, 13, -14, -2, 6, 12, 19, 7, -14, 0, 8, -2, -34, -13, -11, 44, 33, 14, -10, 2, 7, 12, 7, 6, 32, 36, 16, 3, 2, 1, 12, 28, 37, 29, 15, 6, 11, 38, 24, 32, 45, 59, 27, 9, -4},
    '{0, 2, -18, 14, -5, 0, 21, -27, -40, -46, -7, 0, 22, 10, -18, 0, -32, -39, 35, 53, 32, 1, 28, -6, 12, 2, 12, 23, 30, 2, -12, -8, -28, -29, -20, -21, -2, -2, 12, 0, 7, 13, 19, 18, 15, 18, 23, 53, 5, 0, -17, -20, 5, 11, 9, 12, 15, 26, 16, 14, 0, 3, 35, 55, -31, 32, 1, 11, 18, 15, 0, -4, 4, 4, 5, 6, -4, -13, 27, 14, -33, 15, -2, 10, 10, 17, -11, -21, -26, -38, -24, -1, -8, -26, 40, -12, -26, 8, 5, 10, 7, 25, -10, -2, -11, -7, -1, -9, -13, 1, 28, 3, 9, 6, -1, 5, -4, 9, 3, 12, -2, 9, 11, 19, 5, 22, 0, -18, 10, -10, 2, 19, 15, 11, 8, -1, 2, 7, 16, 14, 13, 11, 0, -32, -12, -2, 7, 5, 6, 4, 13, -3, -13, 12, 17, 11, 6, 10, 4, -41, 1, 13, 7, 15, 8, 2, 5, -6, -12, -8, 3, 10, 6, -3, -22, -42, 24, 10, 14, -6, -12, 0, 2, 1, -11, -16, -5, -1, 2, -8, -25, -42, -11, -2, 7, -12, -7, 7, 15, 10, 8, 15, 5, -11, -5, -24, -19, -13, -19, 33, 0, -29, -7, -1, 3, -1, 5, 16, 1, -1, 0, -9, 0, 6, 27, 30, -4, 7, 18, 19, 21, 15, 21, 27, 20, 17, 22, 20, -32, -31, 4, 24, 50, 45, 31, 6, 20, 37, 15, 46, 44, 8, 50, 47, 7, 0},
    '{-1, 1, -4, -24, -16, -33, -55, -31, -10, -4, -35, -40, -71, -50, -11, 4, 24, 5, -16, -2, 22, 0, -7, -8, -6, -9, -22, -7, -32, -29, -5, -25, 27, 35, -3, 1, 11, 11, 20, 5, 9, 11, 1, 6, 0, -8, 2, -3, 0, 1, 3, 9, 11, 3, 3, 0, 4, 7, -4, 8, 0, 0, 9, 17, 23, 10, 14, 9, 0, 9, 9, 7, 3, 4, 0, 2, 3, 11, 10, 23, -24, -5, -1, -1, -3, 1, 15, 16, 8, 7, 8, 5, 11, 12, 22, 8, -32, 12, 8, -13, -21, -15, 17, 23, 9, 10, 13, -2, -16, -15, -2, 29, -37, -5, -4, -22, -22, -15, 7, 17, 14, 8, 13, 6, -16, -36, -33, -4, 13, -25, -6, -29, -23, -13, -6, 6, 9, 2, 5, 1, -6, 3, 12, 23, 16, 9, 15, -18, -17, -19, -42, -17, -3, -4, 12, 19, 16, 29, 29, -10, -11, 41, 23, 17, 4, -11, -18, -22, -9, 2, 0, 15, 9, -5, 1, -58, -29, 17, 13, 18, 8, 4, -2, -4, -7, -4, -5, 11, 4, 2, -26, -50, -4, 7, -18, -4, 5, -1, 3, 5, -3, -13, -5, 6, 7, 3, -44, 6, 12, 28, -6, -16, -7, 0, 6, 0, -4, -5, 13, 7, -4, 5, -17, -4, -21, 11, 1, 8, 6, 12, 11, 24, 0, 1, 6, 6, -12, 5, -3, -39, -3, -11, -21, -14, -36, -24, -1, -15, -27, 4, 16, 1, -29, -8, 9, -11},
    '{-1, -4, 4, 4, -8, 24, 11, -13, -33, -41, -54, 72, 58, 60, 19, 3, 32, 29, 26, -12, -15, 15, 12, -98, -104, -64, -46, 1, 3, 14, 32, 11, 34, 36, -24, -17, 13, 26, -18, -42, -14, -7, -15, 4, -3, 9, -36, -39, 13, 19, -14, -8, 2, 13, -38, -28, 2, -1, 4, 1, 0, 17, -17, 12, 12, 9, -14, -16, -15, 4, -26, -20, -2, 20, 18, 13, 2, 1, -44, 2, 15, 17, -33, -20, 6, 24, -18, -48, -1, 40, 14, -11, -11, -5, -23, 6, -3, -17, -16, -35, 0, 8, -36, -20, 26, 27, 8, -3, -1, -9, -16, 0, -9, 17, -4, -7, -16, -22, -27, 9, 22, 11, 2, -10, 15, 8, 13, 4, 36, 38, -7, -19, 7, 1, 2, 11, 6, 10, 10, -8, 2, -11, 4, 22, 36, 34, -24, -40, -3, 8, 17, 18, 4, -8, -20, -27, 10, 12, 26, 36, 9, 22, -42, -41, -15, 7, 17, 29, -32, -30, -10, -9, 13, 20, 19, 34, -30, -30, -17, -12, -3, -1, 16, 9, -46, -23, -10, -21, -5, -19, -1, -4, -31, -38, -3, 6, -3, 6, -9, -4, -9, -20, -2, 28, 26, 5, 13, 7, -21, -41, 4, 19, 3, 4, -1, 12, 11, -14, -12, 16, -1, 5, 14, 35, 2, -32, 13, -7, 10, 2, 2, 6, 8, -32, -29, -22, -11, 5, -13, -1, 0, 29, 22, 24, 47, 5, -3, 14, 0, -26, -35, -49, 7, 15, -28, 4},
    '{-4, -3, 32, 15, 13, 4, 41, 17, -6, 24, 6, 8, 15, -9, 18, 3, 23, 35, -2, 14, 23, 1, 23, 68, 57, 38, 3, -15, -10, 18, 20, 11, 40, 24, -18, 9, 21, 16, 19, 33, 40, 35, 22, 4, -4, -21, -33, 22, 0, -34, -16, -18, -10, -5, -3, -6, 0, 11, 21, 26, 15, -17, -25, -27, 45, -21, 3, -3, 3, -17, -13, -23, -4, 32, 40, 27, 15, 3, -10, -7, 47, 11, -11, -37, -29, -31, -26, -26, -4, 22, 14, 25, 17, 27, -3, -10, 23, -3, -44, -29, -8, -4, -7, -11, -5, -18, -13, 19, 24, 7, -25, -31, -5, -19, -2, 3, 12, 19, 6, -5, -17, -27, -6, 10, 12, -9, -37, -43, -1, -20, 18, 1, -5, -5, -3, -2, -2, -7, 5, -5, 5, -7, -19, 8, 13, -18, 10, -5, -12, 1, -5, -8, -1, 4, -10, -24, -14, -9, -10, 37, 12, -20, -8, -12, -1, 6, 4, -3, 4, 9, -12, -25, -17, -13, -19, 25, 3, -9, 2, 14, 9, 5, 18, 13, 12, -1, -12, -22, -16, -10, -5, 35, 65, 60, 1, 7, 7, 6, 5, 5, 2, -2, -5, -23, -30, -14, 32, 34, 37, 37, 0, 2, 3, 4, 12, 18, 11, 12, 21, -28, -14, 15, 35, 14, -23, 18, -14, -6, -1, 6, -9, 8, 0, -6, -11, 17, 11, -24, 10, -1, 2, -6, -42, -35, 14, 19, 8, -4, -23, -19, -37, 4, -10, -34, -4, -4},
    '{-2, -4, -4, 8, 9, -1, 4, 4, 2, 27, 43, 26, 2, 2, -2, 0, 3, 1, 4, -4, 4, -15, 0, -13, -26, -19, 26, 25, 3, -14, -24, -18, -3, 20, 2, 3, -5, 3, 4, 2, 15, 9, 4, -11, 7, 27, 32, 16, 39, 3, 1, -1, 3, 15, -2, -1, 4, 4, 14, 9, 6, 7, 33, 29, 57, -7, 1, 0, 1, 4, -1, 3, 13, 23, 22, 22, 1, -11, 2, 46, -18, 10, 8, 1, 9, 3, 0, 2, -18, -33, -32, -18, -4, -7, -5, 43, -10, 18, -3, -4, -7, -9, -14, -9, -28, -18, -25, -41, -33, -51, -23, 45, 20, -8, -6, -11, -22, -14, -1, 15, 16, 4, 2, -3, -15, -36, -49, -38, 28, -28, -13, 9, 6, 12, 13, 5, -1, -7, -4, 5, -2, -9, 9, 9, 29, 30, -1, -11, 4, 18, 30, 19, 3, -10, 2, -5, -4, 6, 24, 32, 40, 43, -6, -52, -52, -54, -53, -41, -16, -7, -3, 8, 0, -5, 22, -5, 44, 43, 5, -30, -32, -44, -28, -11, 6, 14, 8, 15, 2, 0, 43, 32, 17, 32, 27, 2, 9, 6, 31, 19, 7, 5, -2, 16, 0, -12, 6, 15, 22, 55, 51, 22, 14, 12, 18, 1, -1, -1, -7, -3, -5, -25, -10, -5, -18, 27, 33, 40, 35, 34, 23, 16, -3, 8, 11, 4, 29, 5, -4, -9, -2, 11, 27, 15, 0, 16, 19, 8, 7, 17, 3, 12, 22, 32, 23, 0},
    '{-3, -5, -30, -3, 3, 33, 8, -9, 8, -14, 12, 14, 2, -3, 16, 1, 0, -30, -28, 7, 30, 10, 26, -10, -13, -26, -11, 7, -13, -3, 23, 17, 0, -6, 19, 27, 35, 15, 20, 14, -13, -17, -22, -11, 8, 12, 26, 22, 25, 37, 31, 32, 22, 9, 0, 4, -4, 6, -15, -12, -7, 10, 21, 15, 4, 50, 22, 3, -1, -4, 5, 7, -5, -10, -5, -3, 5, 4, 12, 27, 12, 7, -3, -11, -1, -6, -8, -3, -12, -13, -6, 11, 32, 25, 17, 48, -31, -3, -22, -5, 15, -15, -23, -24, -20, -15, -11, 4, 6, -1, 8, 33, -30, -11, -21, -8, 1, -18, -10, 10, 12, -4, -4, 2, -1, -21, 19, 49, 40, 21, -1, 14, 7, -3, 15, 30, 25, 5, 23, 29, 5, -5, 3, 59, 45, 32, 22, 17, 11, -4, -3, 20, 18, 15, 23, 25, 16, 16, 18, 52, 21, 37, 24, 4, -5, -24, -23, 5, 6, 14, 7, -4, 7, 7, 27, 44, -25, 12, 0, -5, -14, -19, -14, -3, 8, 8, -13, -15, -8, -13, -39, -8, -23, -11, -14, -17, -6, -13, -3, 4, 2, -2, -27, -13, -12, -6, -36, -32, 25, -23, 1, 3, 8, 0, 5, -1, 4, 2, -19, -13, -13, -13, -13, -15, 13, 25, 28, 7, -13, -3, 10, -1, 3, 1, -25, -34, -34, -41, -42, 17, 4, 9, -40, -37, -20, 24, 12, -9, 1, -2, 3, -10, -31, -41, -52, 11},
    '{3, -4, -30, -22, -19, -12, 3, 17, -6, -60, -53, -26, -7, 4, -7, 2, -1, -29, -3, -11, -5, -23, -5, -25, -18, -43, -35, -8, -17, -31, -34, -22, -23, -32, 3, -7, -6, 1, 2, 0, -4, -4, 4, 22, 15, 17, 0, -17, 14, -18, -5, 5, -4, -6, -17, -11, -16, -13, 1, 14, 23, 44, -6, -20, 0, 15, 12, 6, -13, -14, -18, -12, -15, -6, 13, 11, 14, 16, -9, -9, 0, 4, 16, -13, -7, -5, -12, -3, -5, 13, 16, 2, -8, -25, -11, -12, 12, -4, -9, -19, -6, 6, 15, 20, -9, 16, 7, -19, -30, -51, -38, -54, 9, -18, -15, -14, 4, 3, 19, 5, -14, 9, 2, -11, -6, -37, -51, -58, 18, 13, 2, -15, 10, 16, 9, -10, -16, 9, 9, 13, 12, -9, -27, -18, 10, 8, -6, -7, 18, 23, 16, 8, -3, 11, 17, 14, -1, -2, -12, -21, -11, 12, -10, -12, 9, 11, 10, 11, 12, 6, 12, 9, -2, -13, -21, -44, 5, 7, -2, -5, -7, -11, -8, -6, 2, 14, 11, -3, -11, -32, -39, -20, 9, 0, -15, -17, -28, -19, -8, -5, 4, 9, 12, 4, 7, -7, -37, -13, -9, -16, -26, -14, -4, 5, 8, 2, 11, 12, 22, 14, 1, -15, -31, 13, 9, 11, -24, -23, -17, 4, 2, -5, 4, 4, 5, -15, -7, -1, -30, -14, 2, 11, -3, -1, -15, -20, -31, -21, -14, -3, -8, -42, -25, -16, -37, -14},
    '{-4, -3, 0, 25, 12, 23, 47, 47, 33, 28, 28, 11, -5, -20, 6, -2, 22, 25, -30, 16, 25, 34, 56, 62, 35, 9, -3, -23, -12, 35, 19, -19, 32, 8, -23, 8, 29, 16, 31, 29, 25, 20, 16, 2, -1, -18, -10, 30, -29, -24, 0, 4, -5, -22, -16, 5, 24, 32, 27, 16, 8, -19, 5, 5, -30, -17, 15, 2, -9, -20, -23, -6, 15, 29, 29, 23, 20, 10, 3, 3, 6, 15, 1, -13, -8, -3, -5, -12, -15, 3, 1, 13, 10, 32, 25, 22, -7, 3, -31, -25, -9, -11, 2, -11, -4, -2, 3, 14, 20, 21, 1, -6, -20, -10, -19, -21, -6, 3, -12, -4, 17, 3, -4, -3, -1, -11, -30, -25, -8, -27, -8, -12, -13, -8, -3, 3, 12, -9, -17, -22, 1, 1, -5, 31, 17, -8, 3, 7, 4, 7, 1, -12, -17, -10, -16, -25, -1, 9, -3, 32, 7, -11, -18, 4, 5, -1, -25, -39, -14, 1, -5, -14, -22, -7, -19, 8, -2, -12, -8, 6, -3, -11, -15, -6, 7, 11, 12, 1, -19, 10, -14, -6, 44, 39, -6, 9, 15, 16, 22, 17, 15, -6, -7, 7, -10, -6, 2, 20, 11, 25, -9, -4, 13, 21, 24, 17, 7, 11, 12, 15, 9, 16, 24, -11, -16, -4, -28, 2, 21, 22, 14, 18, 8, 26, 20, 20, 8, -15, -9, -12, 2, 2, -18, -6, 16, 32, 36, 21, 27, -7, -9, -14, -9, -43, -4, -1},
    '{-4, -1, -28, -8, -23, -39, -24, 22, 21, -31, -20, 8, -17, -27, -19, 3, -21, -29, 16, -25, -49, -38, -27, -13, -6, -14, 15, 20, -4, -28, -24, -24, -38, -3, 41, 13, -45, -40, -21, -1, 4, 5, 8, 1, -3, 11, 16, -3, 18, 38, 25, 12, -17, -28, 7, 15, 15, 7, 12, 11, 1, -1, 12, 23, -30, 37, -21, -32, -29, -26, 13, 24, 10, 10, 16, 7, 8, 8, 31, 30, -40, -25, -52, -44, -39, -30, 27, 25, 10, -6, -4, -10, 1, -2, 52, 5, -20, -1, -9, -33, -61, -29, 21, 15, -10, -6, 7, 3, -12, -3, 27, 23, -7, 2, -24, -32, -28, -1, 16, 4, 7, 5, -11, 1, -16, -25, 3, -9, -7, -26, -3, -19, -8, 2, -5, 0, 13, 16, -9, -11, 0, -9, 19, -27, -51, -20, 13, 5, -2, -10, -7, 4, 11, 21, 10, -19, -17, -10, -29, -61, 0, -19, -8, 1, 2, 3, -5, 3, 16, 19, 3, -17, -30, -19, -2, -24, 26, -38, -17, -18, -8, 2, -1, 6, 8, 6, -5, -26, -46, -35, -12, -28, -37, -45, -8, -3, -3, 4, 17, 20, 3, -8, -17, -44, -67, -55, -9, -47, -37, -23, 15, 8, 5, -7, 11, 20, 11, -11, -43, -55, -53, -15, -22, -43, 16, -20, -3, -1, 7, -1, 19, 21, 7, 5, -47, -51, -27, 33, -23, -27, 4, -2, 25, 15, -2, -23, -19, 11, 4, 33, 51, 2, 8, 56, 1, -4},
    '{-2, -3, -23, -14, -10, -23, 15, 18, 6, -34, -13, 15, 25, 0, 1, -1, -25, -37, -31, -42, -44, -25, -24, -30, -2, -24, -34, -25, -10, -1, -1, -15, -20, -38, -17, -22, -3, 16, 4, -3, 4, 4, 2, 2, 6, 16, 18, 4, -12, 1, 2, -11, 11, 19, -1, 5, 10, 7, 5, -8, 6, 3, -6, -25, -23, 21, 12, -13, -9, -5, -16, 1, 2, 2, 0, 1, 9, -3, 0, -7, 8, 6, -14, 0, -7, -10, -6, 0, 10, -1, -6, 5, 2, -21, -18, 4, 17, -10, -36, -9, -10, -2, 14, 21, 7, 7, -6, 3, 4, -31, -39, -2, 13, -20, -51, -37, -4, 8, 20, 14, 12, 15, 8, 1, 8, -16, -28, -24, -6, -17, -33, -46, -2, 10, 17, 7, 1, 16, 25, 9, 6, -8, -13, -15, 16, -4, -10, -31, 7, 17, 15, 9, 0, 14, 11, -7, -24, 9, -2, -11, 11, 15, -6, -19, 1, 3, -2, 13, 3, -5, -2, -10, -21, 11, 6, 8, 10, 15, -5, -7, -9, -11, -14, -5, -8, -15, -14, -5, -14, -23, -27, 1, 16, -7, -11, -1, -3, -2, 0, 11, -3, -6, -14, -5, -4, -28, -37, 12, -24, -33, -23, -6, 4, 3, 3, 3, 0, -4, 4, 10, 7, -2, -11, 6, 34, -17, 26, 15, -5, -3, 6, -13, -11, -6, -6, -16, -15, 1, -21, -9, 1, -12, 43, 41, 4, -2, -11, -6, -14, -11, 0, -24, -18, -16, -31, -7},
    '{-1, 2, -1, 2, -7, -11, 9, 18, 12, 12, 1, 15, -6, -1, -4, -4, 27, 22, 15, 34, 2, -26, 4, 10, 16, 8, 30, 21, 5, -11, -16, -10, 33, 30, 16, 20, 5, -16, 6, 6, 8, 8, 0, -9, -12, -15, -26, -43, -23, 6, -12, -15, -5, -5, -4, 0, -7, -3, 0, -8, -17, 3, -12, -25, -46, -18, -26, -23, 4, 12, 3, 3, -3, 4, 6, 7, -9, -2, 14, -9, -30, -6, -29, -9, 17, 13, 13, 0, 8, -6, -4, -2, -6, -3, 32, -25, 2, -16, -24, -21, 10, 14, -3, 1, 4, 1, 0, 12, 13, 37, 10, -17, -5, -38, -45, -22, 6, 13, 8, 16, 18, 11, 7, 19, 20, -6, -30, -31, -6, -26, -28, -54, -30, -9, 14, 41, 31, 7, 4, 1, -4, -26, -35, -46, 8, 15, -10, -65, -68, -48, -12, 20, 17, -8, -16, -10, 3, -8, -21, 2, -39, 27, 21, -5, -42, -54, -48, -27, 1, -12, -39, -28, -21, -22, 0, 42, -47, -14, 31, 21, 0, -9, -27, -29, -5, 5, 1, -10, -22, -20, 0, 27, -30, -28, 24, 38, 33, 23, 4, -11, -4, 2, -4, -12, -17, -19, 17, -4, -40, -25, 1, 1, 6, 9, 0, -1, -2, -11, -5, -12, -20, 1, 21, 22, -9, -13, 6, -9, -9, 6, -11, -24, -5, -4, -8, -22, -1, 41, 28, 36, 1, 15, 44, 27, -29, -3, -5, -14, 12, 28, 37, -9, -7, 29, 10, -5},
    '{-2, -2, -12, 21, 34, 50, 25, 0, -18, 6, 6, 2, 30, 19, 18, 4, -24, -16, -39, -11, 10, 26, 36, 13, 22, 12, -13, -24, -1, 22, -1, -19, -24, -22, -2, 17, 17, 19, 0, -3, 1, 15, 5, 2, 9, 2, 11, 22, -19, -1, 25, 10, 5, 2, -10, -7, -5, 11, 1, -3, 4, 9, 5, -1, 26, 12, 41, 9, 3, 6, -6, -7, -4, 1, 2, -8, -2, 14, 2, 22, 15, 23, 14, -1, -5, -4, -21, -6, 3, 13, 11, 13, 18, 31, -17, -6, -16, 6, 2, -8, -5, -17, -13, 0, -1, -7, -9, -4, 2, 9, -1, -19, -19, 8, -11, -13, -9, -2, 9, 21, -8, -9, -9, -7, 1, 0, 16, 13, 12, 29, -2, -5, -1, 11, 14, 22, 9, 2, 0, -10, 0, 6, 22, 57, 44, 28, 3, -3, 8, 15, 12, 17, 13, 10, 0, 12, 19, 18, 35, 53, -26, -4, 11, -8, -5, -1, -1, 5, -5, 10, -5, 0, 8, 7, 9, 23, -33, 15, -5, -6, 9, 0, 5, 5, 12, 4, -8, -10, 7, 0, -14, 38, 44, 62, -2, 7, 19, 5, 15, 8, 2, -8, -12, -1, 4, 7, -26, 11, 40, 33, 3, 12, 14, 16, 19, 26, 8, -1, -6, -1, 7, -2, -30, -24, -6, -1, -22, -4, -25, -16, -2, 5, 8, -1, -7, -29, -27, -27, -18, -2, -3, -38, -44, -34, -27, -34, -14, -39, -65, -26, -4, -50, -60, -36, -23, 8},
    '{-2, 1, 14, -29, -14, 17, -12, 0, -2, 21, 13, 0, -19, -13, 21, 4, -22, 3, -12, -27, -46, -7, -1, 4, -9, -8, -25, -7, 20, 4, 38, 40, -24, -11, -13, -41, -43, -27, -23, -33, -26, -14, -7, -12, -1, -9, -5, -10, 7, 27, 11, -5, -10, -9, -34, -21, -9, -6, -4, -19, -2, -9, -10, -1, 59, 13, -3, 8, 6, 1, -7, -7, -14, -7, -5, -4, 7, 8, 5, -10, 55, 9, 1, 0, -13, -15, 7, 17, 8, 1, 3, 5, -6, 2, 3, -6, 66, 7, -27, -18, -16, -18, 25, 35, 6, -4, 7, 12, -16, -31, -26, -33, 50, 3, -19, -10, 6, 10, 42, 24, -7, 1, 21, 2, -21, -10, 1, -1, 33, 35, 16, 19, 8, 13, 28, 3, -6, 23, 30, 7, 6, 51, 48, 51, 14, 19, 20, 11, 9, 11, 26, 8, 16, 44, 38, 7, 27, 19, 24, 63, 54, 11, 19, -2, 4, -2, 0, 3, 26, 34, 18, -4, 15, 6, -3, 36, 51, 37, 11, -21, -13, -19, -7, -8, 0, 0, -5, -11, 1, -7, -22, 7, -15, 1, 3, -23, -21, -12, -20, -21, -33, -29, -19, -26, -12, -18, -20, -6, -32, -17, -11, 0, -3, 6, -7, -19, -20, -20, -23, -26, -14, -4, -7, -23, -8, -13, 13, -15, -17, -8, -6, 0, -1, -21, -4, -3, -2, 10, 29, 33, -2, 23, -34, -36, -15, -7, -12, -5, 1, -5, -27, 22, 6, 0, 2, 19},
    '{-3, -5, -32, -31, -27, 3, -45, -17, 19, -15, -42, -47, -68, -41, 7, 1, 21, -25, 3, 13, 0, 5, 9, -17, -30, -19, -7, -6, -19, -30, 5, 7, 7, 17, 11, -8, -35, 3, 32, 13, 1, 4, 1, 2, -5, -1, 18, -24, 1, 24, -25, -49, -41, -12, -2, -10, 9, 19, 15, 6, 4, 1, 26, 14, -45, -40, -55, -51, -23, -16, 1, 12, 24, 3, -11, 0, -6, -10, 22, 19, -52, -40, -17, -18, -12, 1, 18, -2, -18, -25, -8, -15, -10, -17, -4, -9, -47, 1, 12, -1, -18, -7, -9, -21, 3, -2, -9, 1, -5, -17, -21, -23, -44, -11, -21, -21, -30, -23, -22, 6, 26, 13, -5, 9, 4, -22, -25, 20, -42, 4, -19, -9, -15, -26, -22, -8, 4, 18, -4, 8, -13, -20, 2, 29, -19, 39, 7, 13, -2, 0, -13, 2, 14, 19, 11, 9, -6, -6, 7, 17, -22, 33, 11, 36, 33, 30, 3, 4, 27, 13, 3, 3, -8, -5, 0, 6, -26, 1, 15, 9, 0, 19, 0, 2, 12, 13, 6, 10, 3, 31, 52, 8, -13, 7, 12, -4, -16, -6, -12, -7, -8, 8, 9, 12, -2, 32, 65, -19, 17, 25, 4, -30, -25, -20, -2, -18, -15, 3, -7, 9, 6, 52, 76, 29, 11, 20, -26, -12, 0, 7, 0, -1, 5, 23, 13, 27, 29, 25, 36, 12, 4, 9, 11, 5, 8, 30, 30, 27, 48, 34, -15, -12, 34, 43, 32, 6},
    '{-1, 2, 32, 29, 21, 24, 64, 38, 9, 21, 4, 19, 25, 25, -7, 2, -6, 36, 46, 33, 8, 17, 39, 39, 52, 9, -37, -21, -18, -1, 5, 0, -8, 8, 7, -10, -12, 0, 6, 25, 27, -3, -35, -48, -27, -15, -16, -24, 13, 2, 21, 3, -9, -15, -14, -11, -32, -27, -18, -8, -11, -3, -10, 1, 58, 15, 28, 20, 18, 22, 12, -14, -41, -18, -6, -22, -4, 14, 30, 9, 73, 20, 29, -1, 11, 18, 34, 2, -21, 20, 15, 9, 27, 20, 31, -3, 57, 18, 8, -10, -7, 13, 23, -15, -17, 28, 22, 13, 15, -1, 19, 10, 38, 15, -10, -2, 1, 12, 14, -30, -22, 0, 6, 6, 8, 9, 35, -2, 70, 32, 12, 17, 14, 12, 8, -9, 0, -11, -11, -5, 0, 26, 5, -47, 31, 16, -3, -1, 4, 7, -4, -4, 13, -14, -2, 6, 9, 0, -9, -46, 26, -37, 13, -9, -14, -4, -17, 0, 6, -4, 7, -7, 6, 12, 13, 4, 39, -16, -18, -1, -1, -9, -2, 3, 1, -10, -9, -15, -17, -13, -22, -10, -2, -1, -44, -10, 8, 12, -4, 2, -3, -3, -7, -14, -10, -3, -5, 38, 5, -3, -20, 5, -4, 9, -2, 14, 8, 6, -9, -21, -12, -8, -10, 32, -11, 18, -4, -8, -17, -19, -9, -4, 4, 7, -3, -26, 0, 15, 11, 3, -2, -2, -49, -39, -25, -28, -22, -26, -32, -23, -25, -17, -23, 5, 1, -1},
    '{-2, -3, 5, 31, 36, 48, 27, 23, 64, 84, 76, 66, 42, 21, 11, 0, 19, 28, 22, 20, -4, 20, -25, -37, -38, -8, -3, -1, 1, 37, 11, 2, 27, 11, -2, -11, -2, 1, -31, -31, -18, 8, 18, -2, -19, 2, 18, 42, -35, -24, -14, -17, 3, -7, -2, 8, 6, 9, 3, -3, 1, 9, 23, 6, -14, -17, 2, 1, 10, -2, 6, 8, -2, -7, -2, 2, 3, 4, -25, 1, 15, -9, 10, 8, -2, 2, 2, 4, -5, -18, -20, -14, -21, 4, -20, 23, 19, -22, 8, 6, 4, 0, 9, -15, -6, 7, -15, -19, -8, -2, -18, -18, 24, 18, 3, 0, 5, 2, -22, -30, -15, -10, -3, -3, 12, -11, -12, 13, -21, 7, -11, 6, -5, -10, -36, -11, -2, -20, -1, 4, 5, -17, -11, 30, -27, 6, -5, 7, -25, -46, -37, 12, 26, 12, -4, 1, -11, 1, 27, 30, 1, 0, -14, -29, -31, -47, -16, 30, 29, 12, 4, 3, -7, -5, 22, 31, 31, 12, -11, -20, -20, -11, 25, 30, 25, 13, 16, 5, -8, -6, 29, 69, 5, 17, 5, -10, -11, 9, 19, 16, 21, 24, 16, -2, -3, 16, 35, 36, 19, -13, 4, -17, -5, 7, 0, 10, 17, 11, -3, 9, 25, 41, 1, 0, 7, -27, -47, -39, -28, -45, -20, -12, 14, 5, 15, 10, 15, 36, 45, -4, 2, -7, -19, -10, 18, -38, -27, -4, 18, -28, -9, 21, 3, -4, 12, 1},
    '{0, 1, 14, -2, 4, -14, -15, 12, 21, 19, 55, 73, 51, 41, 15, 4, 3, 8, -15, -23, -25, -12, 12, 10, -32, -22, 22, 4, -23, -3, 36, 31, 21, 21, -47, -21, -13, -21, -18, -30, -22, -24, -5, -14, 6, 15, -5, 16, 25, 12, -24, -20, -9, -7, 0, 1, 6, -5, 7, 5, 26, 5, 1, -5, 39, 6, -10, -12, -3, -3, 15, 29, 27, 33, 32, 23, 23, 18, -12, -7, 38, -16, 4, -9, -13, 0, 12, 22, 17, 17, 22, 10, 3, 28, 17, -9, 44, -18, -15, 1, -6, 6, 12, -1, -31, -32, -10, -3, -7, -3, 20, 46, 45, -8, -28, -4, 4, 13, 7, -21, -33, -38, -20, -24, -24, -16, 19, 26, 42, -4, -12, 6, -6, 0, 6, -12, -13, -18, -20, -24, -5, 10, 13, -8, -15, -14, -10, -8, 0, 18, 11, -9, -24, -8, -17, -8, 5, 6, -15, -1, -43, -21, -11, -12, -3, 9, -6, -13, -13, -7, -9, 0, 4, -13, -47, -7, 17, 1, 8, 13, 14, 9, -5, -6, -6, -3, -7, -2, -5, -25, -39, 26, 28, 17, 16, 11, 5, 14, 5, 5, 7, 8, 13, 0, -10, 22, 23, 0, 44, 28, 32, 26, 6, 5, 2, 11, 17, 20, 19, 2, -5, 25, 36, 4, -4, 13, 1, 1, 25, 14, 10, 30, 17, 21, 36, 48, 37, 23, 38, 28, 0, 11, -41, -34, 9, -9, -1, 5, 11, 7, 15, 49, 26, 42, 42, 18},
    '{1, 0, -13, -18, 6, 6, -20, -28, 12, 2, -32, -13, -35, -40, 10, 4, 27, 26, -13, -10, 26, 10, 3, -8, -6, -8, -19, -9, -2, 4, -8, -25, 25, 45, 23, 15, 16, 11, 31, 27, 12, 12, 2, 2, 0, 2, 21, 14, -18, 7, 9, 8, 8, 8, 17, 8, 5, 7, 2, 2, -6, 8, 32, 24, -30, 0, 10, -2, 3, 1, -3, 11, 18, 9, -9, -1, -8, 7, 16, 31, -40, -2, -12, -3, -4, 1, -1, 7, 9, -9, -14, -5, 1, 7, -16, 5, -57, -13, -2, -3, -1, -9, -7, 10, 16, -6, -14, -4, -9, -7, -2, 13, -44, -3, -8, -1, -9, -10, -6, 30, 28, 7, 4, 13, 0, -15, -13, 23, -32, -15, -23, -5, -7, -13, -6, 22, 20, 13, 3, -3, -12, -20, 0, 18, 14, 18, 3, -3, 6, -3, -25, 6, 8, 1, 1, -2, -9, 10, 15, -5, -40, 17, 19, 11, 2, -6, -26, -13, -2, 4, 3, 10, 1, 10, 5, -17, -34, -5, 5, 14, -4, 2, -25, -23, 1, 12, 10, 18, 14, 9, -3, -24, 26, 30, -1, 10, 10, 4, 3, -6, -1, 0, -3, 14, 6, -1, -23, -19, 19, 40, -1, -11, 2, 3, 2, -5, -13, -3, 3, 16, 11, 8, -5, 1, -14, 0, -27, 0, 7, 16, 11, 0, -4, 0, 3, -4, -1, -20, -19, -26, 0, -6, -6, 5, -2, 12, 23, -8, -1, 12, 17, -27, 8, 6, 5, -6}
};

// 第1层Bias (int32)
logic signed [31:0] layer1_bias [0:63] = '{
    1392, 385, 2325, 1641, -479, 2640, -179, 1308,
    2541, 418, 1414, -1259, 1784, -381, 919, 440,
    52, -1165, -2276, 549, -623, 1069, 259, 1201,
    153, 37, -338, 1365, -847, 1026, -366, 994,
    251, 1590, 867, 137, 146, 1038, 2526, 565,
    1328, 481, 1948, 297, -1076, -387, 1646, 847,
    64, -90, -176, 2549, -187, -16, 2347, -401,
    1498, 1490, 1535, 1406, 1439, 147, 222, -112
};

// 合并的Scale参数
logic [31:0] merged_scale = 32'b00111010100101110011110001110101;

// 前16个输入 (int8)
logic signed [7:0] input_16 [0:15][0:255] = '{
    '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 10, 8, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 85, 79, 57, 43, 42, 42, 42, 36, 10, 0, 0, 0, 0, 0, 0, 25, 49, 56, 82, 88, 93, 94, 92, 109, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 5, 8, 9, 52, 96, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 98, 60, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 55, 96, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 89, 50, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 65, 92, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 104, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 90, 71, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 64, 112, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 104, 96, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 49, 25, 1, 0, 0, 0, 0, 0, 0, 0},
    '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 18, 30, 29, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 69, 109, 114, 115, 77, 5, 0, 0, 0, 0, 0, 0, 0, 0, 2, 52, 113, 69, 41, 74, 105, 16, 0, 0, 0, 0, 0, 0, 0, 0, 2, 42, 56, 6, 10, 84, 99, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 48, 113, 71, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 98, 96, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 83, 108, 36, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 37, 115, 70, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 89, 107, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 123, 54, 4, 2, 0, 0, 2, 8, 15, 12, 1, 0, 0, 0, 0, 50, 125, 93, 77, 76, 58, 57, 76, 88, 96, 81, 19, 0, 0, 0, 0, 25, 88, 97, 103, 119, 111, 94, 86, 72, 55, 38, 11, 0, 0, 0, 0, 0, 9, 12, 16, 24, 22, 13, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 35, 44, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 66, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 84, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 81, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 71, 71, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 90, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 47, 90, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 73, 65, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 96, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 106, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 67, 90, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 53, 36, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 43, 79, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 24, 98, 122, 56, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 97, 123, 124, 97, 56, 8, 0, 0, 0, 0, 0, 0, 0, 0, 6, 78, 126, 124, 107, 97, 115, 51, 2, 0, 0, 0, 0, 0, 0, 1, 46, 117, 116, 75, 24, 14, 87, 105, 39, 1, 0, 0, 0, 0, 0, 2, 61, 118, 54, 6, 0, 0, 40, 116, 81, 5, 0, 0, 0, 0, 0, 5, 71, 94, 4, 0, 0, 0, 40, 117, 91, 9, 0, 0, 0, 0, 0, 12, 98, 90, 0, 0, 1, 28, 94, 119, 62, 2, 0, 0, 0, 0, 0, 13, 102, 92, 10, 23, 46, 103, 125, 89, 14, 0, 0, 0, 0, 0, 0, 9, 85, 115, 93, 117, 122, 123, 110, 39, 0, 0, 0, 0, 0, 0, 0, 2, 40, 102, 124, 124, 121, 87, 31, 5, 0, 0, 0, 0, 0, 0, 0, 0, 3, 21, 67, 74, 46, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 13, 1, 0, 0, 1, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 70, 4, 0, 0, 10, 46, 7, 0, 0, 0, 0, 0, 0, 0, 1, 39, 77, 4, 0, 0, 11, 73, 17, 0, 0, 0, 0, 0, 0, 0, 17, 85, 33, 1, 0, 0, 20, 95, 20, 0, 0, 0, 0, 0, 0, 5, 63, 76, 2, 0, 0, 1, 58, 92, 13, 0, 0, 0, 0, 0, 0, 15, 92, 36, 0, 0, 0, 13, 98, 54, 2, 0, 0, 0, 0, 0, 0, 18, 90, 24, 2, 2, 3, 33, 108, 33, 0, 0, 0, 0, 0, 0, 0, 9, 77, 84, 57, 58, 69, 96, 109, 20, 0, 0, 0, 0, 0, 0, 0, 0, 13, 45, 57, 54, 38, 88, 102, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 3, 69, 102, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 70, 98, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 78, 54, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 15, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 78, 80, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 113, 70, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 66, 123, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 97, 100, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 114, 68, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 65, 114, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 92, 99, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 114, 65, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 52, 108, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 72, 98, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 57, 80, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 15, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 13, 2, 0, 0, 0, 0, 3, 2, 0, 0, 0, 0, 0, 0, 9, 70, 63, 5, 0, 0, 0, 14, 62, 20, 0, 0, 0, 0, 0, 3, 51, 98, 20, 0, 0, 0, 3, 57, 74, 9, 0, 0, 0, 0, 0, 23, 88, 51, 0, 0, 0, 0, 33, 95, 33, 0, 0, 0, 0, 0, 0, 53, 106, 36, 10, 7, 10, 30, 93, 59, 3, 0, 0, 0, 0, 0, 0, 34, 101, 106, 90, 80, 83, 109, 102, 21, 0, 0, 0, 0, 0, 0, 0, 3, 22, 51, 66, 48, 46, 105, 61, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 41, 94, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 85, 69, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 103, 29, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 60, 103, 41, 32, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 53, 105, 77, 29, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 20, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 20, 47, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 98, 111, 37, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 74, 121, 121, 109, 53, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 98, 47, 53, 111, 111, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 97, 21, 21, 103, 115, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 100, 77, 83, 94, 108, 54, 2, 0, 0, 0, 0, 0, 0, 0, 0, 2, 49, 109, 78, 21, 63, 95, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 18, 9, 0, 14, 96, 53, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 92, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 82, 63, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 88, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 49, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0},
    '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 17, 34, 36, 40, 47, 10, 0, 0, 0, 0, 0, 0, 0, 2, 35, 76, 103, 120, 119, 114, 117, 33, 0, 0, 0, 0, 0, 4, 21, 10, 76, 116, 106, 88, 70, 56, 55, 15, 0, 0, 0, 0, 4, 51, 77, 9, 20, 27, 19, 7, 1, 0, 0, 0, 0, 0, 0, 2, 46, 97, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 94, 69, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 115, 104, 58, 26, 22, 14, 16, 4, 0, 0, 0, 0, 0, 0, 0, 12, 83, 119, 122, 112, 110, 106, 105, 72, 10, 0, 0, 0, 0, 0, 0, 0, 7, 29, 48, 92, 124, 114, 118, 117, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 45, 118, 97, 107, 112, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 86, 118, 111, 58, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 49, 31, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 5, 12, 7, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 14, 47, 72, 94, 78, 50, 22, 0, 0, 0, 0, 0, 0, 0, 10, 48, 96, 105, 81, 78, 100, 114, 86, 14, 0, 0, 0, 0, 0, 11, 74, 114, 70, 23, 3, 28, 60, 101, 116, 28, 0, 0, 0, 0, 0, 28, 108, 100, 53, 56, 59, 81, 112, 119, 81, 9, 0, 0, 0, 0, 0, 10, 58, 94, 99, 99, 114, 126, 120, 72, 17, 0, 0, 0, 0, 0, 0, 0, 1, 13, 17, 33, 101, 119, 58, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 83, 122, 79, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 53, 121, 95, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 101, 111, 39, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 61, 123, 64, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 87, 96, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 32, 32, 1, 0, 0, 0, 0, 0, 0, 0, 0},
    '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 31, 34, 61, 60, 41, 14, 1, 0, 0, 0, 0, 0, 0, 0, 3, 57, 113, 101, 94, 91, 108, 91, 21, 0, 0, 0, 0, 0, 0, 0, 13, 99, 86, 26, 14, 11, 46, 108, 67, 4, 0, 0, 0, 0, 0, 0, 23, 98, 28, 0, 0, 0, 2, 68, 100, 15, 0, 0, 0, 0, 0, 2, 55, 90, 8, 0, 0, 0, 0, 39, 104, 21, 0, 0, 0, 0, 0, 11, 86, 50, 0, 0, 0, 0, 0, 35, 103, 21, 0, 0, 0, 0, 0, 15, 89, 22, 0, 0, 0, 0, 0, 36, 103, 21, 0, 0, 0, 0, 0, 34, 99, 20, 0, 0, 0, 0, 1, 57, 101, 17, 0, 0, 0, 0, 0, 37, 100, 20, 0, 0, 0, 0, 31, 97, 61, 2, 0, 0, 0, 0, 0, 20, 94, 33, 11, 11, 18, 49, 96, 79, 14, 0, 0, 0, 0, 0, 0, 9, 81, 100, 94, 94, 100, 114, 90, 26, 0, 0, 0, 0, 0, 0, 0, 1, 17, 73, 91, 91, 80, 47, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 26, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 98, 71, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 68, 74, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 83, 41, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 32, 104, 23, 0, 1, 20, 46, 55, 33, 3, 0, 0, 0, 0, 0, 1, 54, 83, 4, 12, 56, 105, 98, 92, 104, 27, 0, 0, 0, 0, 0, 8, 81, 59, 12, 79, 103, 57, 14, 14, 84, 37, 0, 0, 0, 0, 0, 11, 92, 54, 44, 101, 41, 4, 0, 9, 73, 23, 0, 0, 0, 0, 0, 12, 94, 54, 57, 96, 21, 0, 0, 30, 84, 14, 0, 0, 0, 0, 0, 16, 98, 58, 9, 66, 73, 19, 43, 87, 46, 1, 0, 0, 0, 0, 0, 6, 64, 93, 41, 36, 64, 82, 92, 43, 5, 0, 0, 0, 0, 0, 0, 0, 10, 64, 92, 95, 92, 76, 24, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 15, 17, 13, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 15, 14, 4, 2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 79, 105, 101, 54, 52, 18, 0, 0, 0, 0, 0, 0, 0, 0, 16, 92, 95, 50, 46, 73, 99, 26, 0, 0, 0, 0, 0, 0, 0, 9, 76, 86, 20, 1, 12, 97, 66, 4, 0, 0, 0, 0, 0, 0, 0, 38, 115, 39, 1, 6, 58, 107, 27, 0, 0, 0, 0, 0, 0, 0, 0, 39, 116, 65, 45, 66, 112, 88, 7, 0, 0, 0, 0, 0, 0, 0, 0, 10, 69, 101, 98, 81, 101, 51, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 14, 12, 50, 109, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 78, 77, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 106, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 47, 102, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 52, 85, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 31, 3, 0, 0, 0, 0, 0, 0},
    '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 18, 23, 12, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 39, 80, 105, 116, 92, 25, 0, 0, 0, 0, 0, 0, 0, 0, 1, 27, 107, 119, 85, 97, 123, 52, 0, 0, 0, 0, 0, 0, 0, 0, 12, 84, 120, 60, 11, 19, 90, 95, 21, 0, 0, 0, 0, 0, 0, 0, 35, 117, 86, 10, 0, 0, 30, 108, 59, 0, 0, 0, 0, 0, 0, 3, 62, 117, 41, 1, 0, 0, 12, 94, 70, 2, 0, 0, 0, 0, 0, 7, 80, 98, 8, 0, 0, 0, 11, 95, 85, 6, 0, 0, 0, 0, 0, 11, 92, 90, 0, 0, 0, 0, 11, 95, 85, 6, 0, 0, 0, 0, 0, 10, 87, 94, 4, 0, 0, 0, 18, 100, 47, 1, 0, 0, 0, 0, 0, 1, 38, 105, 38, 1, 0, 1, 51, 89, 13, 0, 0, 0, 0, 0, 0, 0, 7, 66, 79, 17, 7, 32, 96, 49, 2, 0, 0, 0, 0, 0, 0, 0, 0, 9, 62, 78, 73, 92, 68, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 19, 27, 16, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 77, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 67, 121, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 73, 122, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 59, 120, 52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 74, 125, 59, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 74, 124, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 74, 122, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 74, 122, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 63, 121, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 78, 123, 59, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 111, 105, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 65, 21, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
    '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 15, 24, 52, 82, 81, 56, 23, 1, 0, 0, 0, 0, 0, 0, 0, 37, 99, 90, 76, 62, 33, 8, 2, 0, 0, 0, 0, 0, 0, 0, 0, 27, 104, 43, 7, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 72, 51, 8, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 91, 99, 85, 80, 45, 10, 0, 0, 0, 0, 0, 0, 0, 0, 2, 49, 79, 35, 27, 44, 74, 76, 38, 4, 0, 0, 0, 0, 0, 0, 0, 8, 9, 0, 0, 1, 7, 36, 77, 47, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 80, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 43, 82, 0, 0, 0, 0, 0, 0, 19, 24, 0, 0, 0, 2, 7, 22, 73, 50, 0, 0, 0, 0, 0, 4, 62, 83, 37, 37, 43, 59, 74, 79, 52, 8, 0, 0, 0, 0, 0, 1, 23, 60, 73, 76, 67, 54, 35, 17, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0}
};
